--
-- (C) 2018, ZPUROMGEN, Yosel de Jesus Balibrea Lastre.
--           Automatically Generated ROM file
--           Please do NOT CHANGE!
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity prog_mem is
generic
(
maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
);
port (
		clk : in std_logic;
		areset : in std_logic := '0';
		from_zpu : in ZPU_ToROM;
		to_zpu : out ZPU_FromROM
		);
end prog_mem;

architecture rtl of prog_mem is

	type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

	shared variable ram : ram_type := (
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080e7c0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff2",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"8080e3ce",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c32d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870892a",
   171 => x"70810651",
   172 => x"515170f3",
   173 => x"3871c00c",
   174 => x"7183ffe0",
   175 => x"800c0288",
   176 => x"050d0402",
   177 => x"e8050d80",
   178 => x"78575575",
   179 => x"70840557",
   180 => x"08538054",
   181 => x"72982a73",
   182 => x"882b5452",
   183 => x"71802ea0",
   184 => x"38c00870",
   185 => x"892a7081",
   186 => x"06515151",
   187 => x"70f33871",
   188 => x"c00c8115",
   189 => x"81155555",
   190 => x"837425d8",
   191 => x"3871cc38",
   192 => x"7483ffe0",
   193 => x"800c0298",
   194 => x"050d0402",
   195 => x"fc050dc0",
   196 => x"0870882a",
   197 => x"70810651",
   198 => x"515170f3",
   199 => x"38c00870",
   200 => x"81ff0683",
   201 => x"ffe0800c",
   202 => x"51028405",
   203 => x"0d0402e8",
   204 => x"050d777a",
   205 => x"57548055",
   206 => x"84808086",
   207 => x"8b2d83ff",
   208 => x"e0800881",
   209 => x"ff065372",
   210 => x"882e0981",
   211 => x"06a33880",
   212 => x"7525e538",
   213 => x"75802e8d",
   214 => x"38848080",
   215 => x"e7d05184",
   216 => x"808085c3",
   217 => x"2dff14ff",
   218 => x"16565484",
   219 => x"808086b8",
   220 => x"04728d2e",
   221 => x"b638e013",
   222 => x"527180de",
   223 => x"26ffb938",
   224 => x"75802e92",
   225 => x"38c00870",
   226 => x"892a7081",
   227 => x"06515152",
   228 => x"71f33872",
   229 => x"c00c7274",
   230 => x"70810556",
   231 => x"84808081",
   232 => x"b72d8115",
   233 => x"55848080",
   234 => x"86b80480",
   235 => x"74848080",
   236 => x"81b72d74",
   237 => x"83ffe080",
   238 => x"0c029805",
   239 => x"0d0402d0",
   240 => x"050d8070",
   241 => x"57578177",
   242 => x"54588852",
   243 => x"02a40570",
   244 => x"52598480",
   245 => x"8086ae2d",
   246 => x"76557419",
   247 => x"70848080",
   248 => x"80f52d89",
   249 => x"0bd01227",
   250 => x"78058118",
   251 => x"58585154",
   252 => x"877525e6",
   253 => x"38807625",
   254 => x"a63802a3",
   255 => x"05557515",
   256 => x"70848080",
   257 => x"80f52dd0",
   258 => x"117a2979",
   259 => x"057a8829",
   260 => x"7b1005ff",
   261 => x"1a5a5b59",
   262 => x"51547580",
   263 => x"24e03876",
   264 => x"83ffe080",
   265 => x"0c02b005",
   266 => x"0d0402f4",
   267 => x"050dd452",
   268 => x"81ff720c",
   269 => x"71085381",
   270 => x"ff720c72",
   271 => x"882b83fe",
   272 => x"80067208",
   273 => x"7081ff06",
   274 => x"51525381",
   275 => x"ff720c72",
   276 => x"7107882b",
   277 => x"72087081",
   278 => x"ff065152",
   279 => x"5381ff72",
   280 => x"0c727107",
   281 => x"882b7208",
   282 => x"7081ff06",
   283 => x"720783ff",
   284 => x"e0800c52",
   285 => x"53028c05",
   286 => x"0d0402f4",
   287 => x"050d7476",
   288 => x"7181ff06",
   289 => x"d40c5353",
   290 => x"83fff2e4",
   291 => x"08853871",
   292 => x"892b5271",
   293 => x"982ad40c",
   294 => x"71902a70",
   295 => x"81ff06d4",
   296 => x"0c517188",
   297 => x"2a7081ff",
   298 => x"06d40c51",
   299 => x"7181ff06",
   300 => x"d40c7290",
   301 => x"2a7081ff",
   302 => x"06d40c51",
   303 => x"d4087081",
   304 => x"ff065151",
   305 => x"82b8bf52",
   306 => x"7081ff2e",
   307 => x"09810694",
   308 => x"3881ff0b",
   309 => x"d40cd408",
   310 => x"7081ff06",
   311 => x"ff145451",
   312 => x"5171e538",
   313 => x"7083ffe0",
   314 => x"800c028c",
   315 => x"050d0402",
   316 => x"fc050d81",
   317 => x"c75181ff",
   318 => x"0bd40cff",
   319 => x"11517080",
   320 => x"25f43802",
   321 => x"84050d04",
   322 => x"02f0050d",
   323 => x"84808089",
   324 => x"ef2d819c",
   325 => x"9f538052",
   326 => x"87fc80f7",
   327 => x"51848080",
   328 => x"88fa2d83",
   329 => x"ffe08008",
   330 => x"5483ffe0",
   331 => x"8008812e",
   332 => x"098106ae",
   333 => x"3881ff0b",
   334 => x"d40c820a",
   335 => x"52849c80",
   336 => x"e9518480",
   337 => x"8088fa2d",
   338 => x"83ffe080",
   339 => x"088e3881",
   340 => x"ff0bd40c",
   341 => x"73538480",
   342 => x"808ae904",
   343 => x"84808089",
   344 => x"ef2dff13",
   345 => x"5372ffae",
   346 => x"387283ff",
   347 => x"e0800c02",
   348 => x"90050d04",
   349 => x"02f4050d",
   350 => x"81ff0bd4",
   351 => x"0c935380",
   352 => x"5287fc80",
   353 => x"c1518480",
   354 => x"8088fa2d",
   355 => x"83ffe080",
   356 => x"088e3881",
   357 => x"ff0bd40c",
   358 => x"81538480",
   359 => x"808bac04",
   360 => x"84808089",
   361 => x"ef2dff13",
   362 => x"5372d438",
   363 => x"7283ffe0",
   364 => x"800c028c",
   365 => x"050d0402",
   366 => x"f0050d84",
   367 => x"808089ef",
   368 => x"2d83aa52",
   369 => x"849c80c8",
   370 => x"51848080",
   371 => x"88fa2d83",
   372 => x"ffe08008",
   373 => x"812e0981",
   374 => x"06a93884",
   375 => x"808088aa",
   376 => x"2d83ffe0",
   377 => x"800883ff",
   378 => x"ff065372",
   379 => x"83aa2ebb",
   380 => x"3883ffe0",
   381 => x"80085284",
   382 => x"8080e7d4",
   383 => x"51848080",
   384 => x"82e32d84",
   385 => x"80808af4",
   386 => x"2d848080",
   387 => x"8ca30481",
   388 => x"54848080",
   389 => x"8dac0484",
   390 => x"8080e7ec",
   391 => x"51848080",
   392 => x"82e32d80",
   393 => x"54848080",
   394 => x"8dac0481",
   395 => x"ff0bd40c",
   396 => x"b1538480",
   397 => x"808a882d",
   398 => x"83ffe080",
   399 => x"08802e80",
   400 => x"dc388052",
   401 => x"87fc80fa",
   402 => x"51848080",
   403 => x"88fa2d83",
   404 => x"ffe08008",
   405 => x"b63881ff",
   406 => x"0bd40cd4",
   407 => x"085381ff",
   408 => x"0bd40c81",
   409 => x"ff0bd40c",
   410 => x"81ff0bd4",
   411 => x"0c81ff0b",
   412 => x"d40c7286",
   413 => x"2a708106",
   414 => x"83ffe080",
   415 => x"08565153",
   416 => x"72802ea8",
   417 => x"38848080",
   418 => x"8c8f0483",
   419 => x"ffe08008",
   420 => x"52848080",
   421 => x"e8885184",
   422 => x"808082e3",
   423 => x"2d72822e",
   424 => x"fef538ff",
   425 => x"135372ff",
   426 => x"89387254",
   427 => x"7383ffe0",
   428 => x"800c0290",
   429 => x"050d0402",
   430 => x"f4050d81",
   431 => x"0b83fff2",
   432 => x"e40cd008",
   433 => x"708f2a70",
   434 => x"81065151",
   435 => x"5372f338",
   436 => x"72d00c84",
   437 => x"808089ef",
   438 => x"2dd00870",
   439 => x"8f2a7081",
   440 => x"06515153",
   441 => x"72f33881",
   442 => x"0bd00c87",
   443 => x"53805284",
   444 => x"d480c051",
   445 => x"84808088",
   446 => x"fa2d83ff",
   447 => x"e0800881",
   448 => x"2e973872",
   449 => x"822e0981",
   450 => x"06893880",
   451 => x"53848080",
   452 => x"8eda04ff",
   453 => x"135372d5",
   454 => x"38848080",
   455 => x"8bb72d83",
   456 => x"ffe08008",
   457 => x"83fff2e4",
   458 => x"0c83ffe0",
   459 => x"80088e38",
   460 => x"815287fc",
   461 => x"80d05184",
   462 => x"808088fa",
   463 => x"2d81ff0b",
   464 => x"d40cd008",
   465 => x"708f2a70",
   466 => x"81065151",
   467 => x"5372f338",
   468 => x"72d00c81",
   469 => x"ff0bd40c",
   470 => x"81537283",
   471 => x"ffe0800c",
   472 => x"028c050d",
   473 => x"04800b83",
   474 => x"ffe0800c",
   475 => x"0402e005",
   476 => x"0d797b57",
   477 => x"57805881",
   478 => x"ff0bd40c",
   479 => x"d008708f",
   480 => x"2a708106",
   481 => x"51515473",
   482 => x"f3388281",
   483 => x"0bd00c81",
   484 => x"ff0bd40c",
   485 => x"765287fc",
   486 => x"80d15184",
   487 => x"808088fa",
   488 => x"2d80dbc6",
   489 => x"df5583ff",
   490 => x"e0800880",
   491 => x"2e9b3883",
   492 => x"ffe08008",
   493 => x"53765284",
   494 => x"8080e894",
   495 => x"51848080",
   496 => x"82e32d84",
   497 => x"8080909f",
   498 => x"0481ff0b",
   499 => x"d40cd408",
   500 => x"7081ff06",
   501 => x"51547381",
   502 => x"fe2e0981",
   503 => x"06a53880",
   504 => x"ff548480",
   505 => x"8088aa2d",
   506 => x"83ffe080",
   507 => x"08767084",
   508 => x"05580cff",
   509 => x"14547380",
   510 => x"25e83881",
   511 => x"58848080",
   512 => x"908904ff",
   513 => x"155574c1",
   514 => x"3881ff0b",
   515 => x"d40cd008",
   516 => x"708f2a70",
   517 => x"81065151",
   518 => x"5473f338",
   519 => x"73d00c77",
   520 => x"83ffe080",
   521 => x"0c02a005",
   522 => x"0d0402ec",
   523 => x"050d7678",
   524 => x"7a555555",
   525 => x"80732798",
   526 => x"38735274",
   527 => x"51848080",
   528 => x"8eed2d81",
   529 => x"15848015",
   530 => x"ff155555",
   531 => x"5572ea38",
   532 => x"810b83ff",
   533 => x"e0800c02",
   534 => x"94050d04",
   535 => x"02fc050d",
   536 => x"74518071",
   537 => x"278738ff",
   538 => x"115170fb",
   539 => x"38810b83",
   540 => x"ffe0800c",
   541 => x"0284050d",
   542 => x"0402fc05",
   543 => x"0d7270ff",
   544 => x"b40c83ff",
   545 => x"e0800c02",
   546 => x"84050d04",
   547 => x"ffb40883",
   548 => x"ffe0800c",
   549 => x"04c80883",
   550 => x"ffe0800c",
   551 => x"0402ec05",
   552 => x"0d765480",
   553 => x"0b84d415",
   554 => x"0cff0b88",
   555 => x"d8150c80",
   556 => x"0b88dc15",
   557 => x"0c84d814",
   558 => x"55848053",
   559 => x"80527451",
   560 => x"848080e0",
   561 => x"f02d800b",
   562 => x"88e0150c",
   563 => x"84d41408",
   564 => x"88e4150c",
   565 => x"7484d415",
   566 => x"0c029405",
   567 => x"0d0402d8",
   568 => x"050d7b7d",
   569 => x"70565855",
   570 => x"76802e80",
   571 => x"d0388484",
   572 => x"1708802e",
   573 => x"80c538b8",
   574 => x"15085978",
   575 => x"802eb638",
   576 => x"810b8480",
   577 => x"18087094",
   578 => x"18083172",
   579 => x"11a01908",
   580 => x"59575859",
   581 => x"5a747427",
   582 => x"85387476",
   583 => x"315a7953",
   584 => x"76527751",
   585 => x"782d83ff",
   586 => x"e0800854",
   587 => x"83ffe080",
   588 => x"08802e89",
   589 => x"38800b84",
   590 => x"84180c81",
   591 => x"547383ff",
   592 => x"e0800c02",
   593 => x"a8050d04",
   594 => x"02e0050d",
   595 => x"797b5957",
   596 => x"800b84d4",
   597 => x"18085656",
   598 => x"74762e80",
   599 => x"db388480",
   600 => x"15085473",
   601 => x"78268938",
   602 => x"81145473",
   603 => x"7826ae38",
   604 => x"848c1508",
   605 => x"54739638",
   606 => x"75802e8c",
   607 => x"3873848c",
   608 => x"170c8480",
   609 => x"80938d04",
   610 => x"7584d418",
   611 => x"0c74848c",
   612 => x"16085656",
   613 => x"74c83884",
   614 => x"808093b8",
   615 => x"0474802e",
   616 => x"97387784",
   617 => x"80160831",
   618 => x"892b7505",
   619 => x"8488160c",
   620 => x"74548480",
   621 => x"80949a04",
   622 => x"84d41708",
   623 => x"848c170c",
   624 => x"7584d418",
   625 => x"0c848416",
   626 => x"08802e9a",
   627 => x"38755276",
   628 => x"51848080",
   629 => x"91de2d83",
   630 => x"ffe08008",
   631 => x"5483ffe0",
   632 => x"8008802e",
   633 => x"b5387784",
   634 => x"80170c81",
   635 => x"53755284",
   636 => x"80160851",
   637 => x"b4170854",
   638 => x"732d83ff",
   639 => x"e0800893",
   640 => x"38ff0b84",
   641 => x"80170c83",
   642 => x"ffe08008",
   643 => x"54848080",
   644 => x"949a0475",
   645 => x"8488170c",
   646 => x"75547383",
   647 => x"ffe0800c",
   648 => x"02a0050d",
   649 => x"0402f005",
   650 => x"0d7584d4",
   651 => x"11085454",
   652 => x"72802eb1",
   653 => x"38848413",
   654 => x"08802e9e",
   655 => x"38725273",
   656 => x"51848080",
   657 => x"91de2d83",
   658 => x"ffe08008",
   659 => x"8d3883ff",
   660 => x"e0800853",
   661 => x"84808094",
   662 => x"e704848c",
   663 => x"13085384",
   664 => x"808094b0",
   665 => x"04815372",
   666 => x"83ffe080",
   667 => x"0c029005",
   668 => x"0d0402e8",
   669 => x"050d7779",
   670 => x"55567383",
   671 => x"38825473",
   672 => x"882a53b0",
   673 => x"1608802e",
   674 => x"85387387",
   675 => x"2a539416",
   676 => x"08135275",
   677 => x"51848080",
   678 => x"92c82dff",
   679 => x"5583ffe0",
   680 => x"8008802e",
   681 => x"819a3883",
   682 => x"ffe08008",
   683 => x"84880508",
   684 => x"55b01608",
   685 => x"b2387288",
   686 => x"2b747131",
   687 => x"107083ff",
   688 => x"fe061781",
   689 => x"11848080",
   690 => x"80f52d71",
   691 => x"84808080",
   692 => x"f52d7182",
   693 => x"802905fc",
   694 => x"80881153",
   695 => x"58585151",
   696 => x"53848080",
   697 => x"96b70472",
   698 => x"872b7471",
   699 => x"31822b83",
   700 => x"fffc0616",
   701 => x"83118480",
   702 => x"8080f52d",
   703 => x"82128480",
   704 => x"8080f52d",
   705 => x"7181800a",
   706 => x"29718480",
   707 => x"80290581",
   708 => x"14848080",
   709 => x"80f52d70",
   710 => x"82802912",
   711 => x"75848080",
   712 => x"80f52d56",
   713 => x"7505f00a",
   714 => x"06ff8080",
   715 => x"80881153",
   716 => x"55535459",
   717 => x"575553ff",
   718 => x"55877327",
   719 => x"83387355",
   720 => x"7483ffe0",
   721 => x"800c0298",
   722 => x"050d0402",
   723 => x"e0050d79",
   724 => x"7b5856b0",
   725 => x"1608802e",
   726 => x"81ba3898",
   727 => x"16848080",
   728 => x"80e02d9c",
   729 => x"17080552",
   730 => x"75518480",
   731 => x"8092c82d",
   732 => x"83ffe080",
   733 => x"085883ff",
   734 => x"e0800880",
   735 => x"2e819538",
   736 => x"83ffe080",
   737 => x"08848805",
   738 => x"08547683",
   739 => x"ec158480",
   740 => x"8081b72d",
   741 => x"83ffe080",
   742 => x"08848805",
   743 => x"0877882a",
   744 => x"55557383",
   745 => x"ed168480",
   746 => x"8081b72d",
   747 => x"83ffe080",
   748 => x"08848805",
   749 => x"0877902a",
   750 => x"55557383",
   751 => x"ee168480",
   752 => x"8081b72d",
   753 => x"83ffe080",
   754 => x"08848805",
   755 => x"0877982a",
   756 => x"55557383",
   757 => x"ef168480",
   758 => x"8081b72d",
   759 => x"810b83ff",
   760 => x"e0800884",
   761 => x"84050c76",
   762 => x"a4170cb8",
   763 => x"16085473",
   764 => x"802e9538",
   765 => x"815383ff",
   766 => x"e0800852",
   767 => x"83ffe080",
   768 => x"08848005",
   769 => x"0851732d",
   770 => x"ff0b8480",
   771 => x"190c800b",
   772 => x"8484190c",
   773 => x"02a0050d",
   774 => x"0402d005",
   775 => x"0d7d5780",
   776 => x"705956a0",
   777 => x"1708762e",
   778 => x"81ba3894",
   779 => x"17081852",
   780 => x"76518480",
   781 => x"8092c82d",
   782 => x"83ffe080",
   783 => x"08802e81",
   784 => x"a338800b",
   785 => x"b0180883",
   786 => x"ffe08008",
   787 => x"84880508",
   788 => x"5b5b5574",
   789 => x"83ffff06",
   790 => x"5379ad38",
   791 => x"72198111",
   792 => x"84808080",
   793 => x"f52d7184",
   794 => x"808080f5",
   795 => x"2d718280",
   796 => x"29057081",
   797 => x"05097080",
   798 => x"251a821a",
   799 => x"5a5a5152",
   800 => x"55538480",
   801 => x"8099d204",
   802 => x"72198311",
   803 => x"84808080",
   804 => x"f52d8212",
   805 => x"84808080",
   806 => x"f52d7181",
   807 => x"800a2971",
   808 => x"84808029",
   809 => x"05811484",
   810 => x"808080f5",
   811 => x"2d708280",
   812 => x"29127584",
   813 => x"808080f5",
   814 => x"2d710570",
   815 => x"81050970",
   816 => x"72078025",
   817 => x"7e05841e",
   818 => x"5e5e5751",
   819 => x"5253575d",
   820 => x"5d5383ff",
   821 => x"7527fefb",
   822 => x"38811858",
   823 => x"a0170878",
   824 => x"26fec838",
   825 => x"7583ffe0",
   826 => x"800c02b0",
   827 => x"050d0402",
   828 => x"ec050d76",
   829 => x"538054ff",
   830 => x"5272742e",
   831 => x"81963872",
   832 => x"84808080",
   833 => x"f52d5170",
   834 => x"af2e0981",
   835 => x"068c3870",
   836 => x"81145455",
   837 => x"8480809a",
   838 => x"c4048113",
   839 => x"84808080",
   840 => x"f52d5170",
   841 => x"ba2e9638",
   842 => x"82138480",
   843 => x"8080f52d",
   844 => x"51ff5270",
   845 => x"80dc2e09",
   846 => x"810680d8",
   847 => x"3880dc0b",
   848 => x"83145455",
   849 => x"72848080",
   850 => x"80f52d70",
   851 => x"81ff0652",
   852 => x"5270802e",
   853 => x"bc387181",
   854 => x"ff065170",
   855 => x"802ea938",
   856 => x"7181ff06",
   857 => x"81145351",
   858 => x"70752e09",
   859 => x"81068938",
   860 => x"71538480",
   861 => x"809b8804",
   862 => x"71728480",
   863 => x"8080f52d",
   864 => x"53538480",
   865 => x"809ad604",
   866 => x"81145484",
   867 => x"80809ac4",
   868 => x"04ff1452",
   869 => x"7183ffe0",
   870 => x"800c0294",
   871 => x"050d0402",
   872 => x"d0050d7d",
   873 => x"7f616358",
   874 => x"5d5d5380",
   875 => x"70748105",
   876 => x"09707607",
   877 => x"73257074",
   878 => x"7a250751",
   879 => x"51545b58",
   880 => x"ff547178",
   881 => x"2e098106",
   882 => x"81d63872",
   883 => x"84808080",
   884 => x"f52d5271",
   885 => x"af2e0981",
   886 => x"068c3871",
   887 => x"81145457",
   888 => x"8480809c",
   889 => x"90048113",
   890 => x"84808080",
   891 => x"f52d5271",
   892 => x"ba2e9638",
   893 => x"82138480",
   894 => x"8080f52d",
   895 => x"52ff5471",
   896 => x"80dc2e09",
   897 => x"81068198",
   898 => x"3880dc0b",
   899 => x"83145457",
   900 => x"72518480",
   901 => x"80d8f22d",
   902 => x"800b83ff",
   903 => x"e0800825",
   904 => x"80cf38ff",
   905 => x"1583ffe0",
   906 => x"80085559",
   907 => x"72848080",
   908 => x"80f52d70",
   909 => x"81ff0670",
   910 => x"79327081",
   911 => x"05097080",
   912 => x"251e5e51",
   913 => x"54565679",
   914 => x"7c2e0981",
   915 => x"06993874",
   916 => x"772e9438",
   917 => x"7779258f",
   918 => x"387a1852",
   919 => x"75728480",
   920 => x"8081b72d",
   921 => x"81185881",
   922 => x"13ff1555",
   923 => x"5373ffbc",
   924 => x"387a8480",
   925 => x"8080f52d",
   926 => x"5271802e",
   927 => x"95388480",
   928 => x"80eba451",
   929 => x"84808085",
   930 => x"c32d8054",
   931 => x"8480809d",
   932 => x"a0048480",
   933 => x"80eba451",
   934 => x"84808085",
   935 => x"c32dff54",
   936 => x"7383ffe0",
   937 => x"800c02b0",
   938 => x"050d0402",
   939 => x"d8050d7b",
   940 => x"7d7f6173",
   941 => x"555c5c59",
   942 => x"57848080",
   943 => x"99ef2d83",
   944 => x"ffe08008",
   945 => x"83ffe080",
   946 => x"08565683",
   947 => x"ffe08008",
   948 => x"ff2e80f2",
   949 => x"387f5478",
   950 => x"5383ffe0",
   951 => x"80085276",
   952 => x"51848080",
   953 => x"9b9f2dff",
   954 => x"5583ffe0",
   955 => x"800880d6",
   956 => x"38759338",
   957 => x"83ffe080",
   958 => x"08788480",
   959 => x"8081b72d",
   960 => x"8480809e",
   961 => x"c4047651",
   962 => x"848080d8",
   963 => x"f22d83ff",
   964 => x"e0800879",
   965 => x"52558480",
   966 => x"80d8f22d",
   967 => x"7483ffe0",
   968 => x"80083155",
   969 => x"79752583",
   970 => x"38795574",
   971 => x"53765277",
   972 => x"51848080",
   973 => x"ddfd2d74",
   974 => x"18ff0555",
   975 => x"80758480",
   976 => x"8081b72d",
   977 => x"80557483",
   978 => x"ffe0800c",
   979 => x"02a8050d",
   980 => x"0402e005",
   981 => x"0d797bff",
   982 => x"1e565657",
   983 => x"73ff2e80",
   984 => x"d7387684",
   985 => x"808080f5",
   986 => x"2d707684",
   987 => x"808080f5",
   988 => x"2d70ffbf",
   989 => x"14555954",
   990 => x"59537099",
   991 => x"268938a0",
   992 => x"137081ff",
   993 => x"065951ff",
   994 => x"bf125170",
   995 => x"99268938",
   996 => x"a0127081",
   997 => x"ff065751",
   998 => x"77763151",
   999 => x"709c3872",
  1000 => x"802e9538",
  1001 => x"71802e90",
  1002 => x"38811781",
  1003 => x"16ff1656",
  1004 => x"56578480",
  1005 => x"809edc04",
  1006 => x"80517083",
  1007 => x"ffe0800c",
  1008 => x"02a0050d",
  1009 => x"0402ec05",
  1010 => x"0d7654ff",
  1011 => x"74545572",
  1012 => x"84808080",
  1013 => x"f52d7081",
  1014 => x"ff065252",
  1015 => x"70802e9b",
  1016 => x"387181ff",
  1017 => x"065170ae",
  1018 => x"2e098106",
  1019 => x"85387274",
  1020 => x"31558113",
  1021 => x"53848080",
  1022 => x"9fcf0474",
  1023 => x"83ffe080",
  1024 => x"0c029405",
  1025 => x"0d0402ec",
  1026 => x"050d7678",
  1027 => x"707113ff",
  1028 => x"05555555",
  1029 => x"5573802e",
  1030 => x"9e387184",
  1031 => x"808080f5",
  1032 => x"2d5170a0",
  1033 => x"2e098106",
  1034 => x"8e387175",
  1035 => x"31ff13ff",
  1036 => x"16565353",
  1037 => x"73e43872",
  1038 => x"83ffe080",
  1039 => x"0c029405",
  1040 => x"0d0402d4",
  1041 => x"050d7c7e",
  1042 => x"59598079",
  1043 => x"52578480",
  1044 => x"809fc52d",
  1045 => x"83ffe080",
  1046 => x"08785256",
  1047 => x"8480809f",
  1048 => x"c52d83ff",
  1049 => x"e0800876",
  1050 => x"09708105",
  1051 => x"09707207",
  1052 => x"7a255156",
  1053 => x"565a83ff",
  1054 => x"e08008ff",
  1055 => x"2e8c3876",
  1056 => x"5b73772e",
  1057 => x"09810681",
  1058 => x"f73883ff",
  1059 => x"e0800809",
  1060 => x"70810509",
  1061 => x"70720780",
  1062 => x"25515555",
  1063 => x"75ff2e80",
  1064 => x"e238805b",
  1065 => x"737b2e09",
  1066 => x"810681d4",
  1067 => x"3875ff2e",
  1068 => x"80d13875",
  1069 => x"19810583",
  1070 => x"ffe08008",
  1071 => x"19810571",
  1072 => x"53565784",
  1073 => x"8080d8f2",
  1074 => x"2d83ffe0",
  1075 => x"80087552",
  1076 => x"54848080",
  1077 => x"d8f22d73",
  1078 => x"83ffe080",
  1079 => x"082e0981",
  1080 => x"06819d38",
  1081 => x"73537452",
  1082 => x"76518480",
  1083 => x"809ed12d",
  1084 => x"757a5555",
  1085 => x"83ffe080",
  1086 => x"087b2ea3",
  1087 => x"38848080",
  1088 => x"a3800478",
  1089 => x"51848080",
  1090 => x"d8f22d83",
  1091 => x"ffe08008",
  1092 => x"78525584",
  1093 => x"8080d8f2",
  1094 => x"2d83ffe0",
  1095 => x"80085474",
  1096 => x"52785184",
  1097 => x"8080a086",
  1098 => x"2d83ffe0",
  1099 => x"80087453",
  1100 => x"78525584",
  1101 => x"8080a086",
  1102 => x"2d805b74",
  1103 => x"83ffe080",
  1104 => x"082e0981",
  1105 => x"06ba3883",
  1106 => x"ffe08008",
  1107 => x"53775278",
  1108 => x"51848080",
  1109 => x"9ed12d83",
  1110 => x"ffe08008",
  1111 => x"7b2e9338",
  1112 => x"848080eb",
  1113 => x"a4518480",
  1114 => x"8085c32d",
  1115 => x"848080a3",
  1116 => x"80048480",
  1117 => x"80eba451",
  1118 => x"84808085",
  1119 => x"c32d815b",
  1120 => x"7a83ffe0",
  1121 => x"800c02ac",
  1122 => x"050d0402",
  1123 => x"f0050d75",
  1124 => x"5372802e",
  1125 => x"80d73872",
  1126 => x"84808080",
  1127 => x"f52d7081",
  1128 => x"ff065252",
  1129 => x"70802e80",
  1130 => x"c4388113",
  1131 => x"84808080",
  1132 => x"f52d5170",
  1133 => x"af387072",
  1134 => x"81ff0652",
  1135 => x"547080dc",
  1136 => x"2e098106",
  1137 => x"83388154",
  1138 => x"70af3270",
  1139 => x"81050970",
  1140 => x"80257607",
  1141 => x"51515170",
  1142 => x"802e8938",
  1143 => x"81518480",
  1144 => x"80a3ef04",
  1145 => x"81135384",
  1146 => x"8080a397",
  1147 => x"04805170",
  1148 => x"83ffe080",
  1149 => x"0c029005",
  1150 => x"0d0402e8",
  1151 => x"050d7779",
  1152 => x"55558056",
  1153 => x"848080a4",
  1154 => x"b4047181",
  1155 => x"15555371",
  1156 => x"a02ea138",
  1157 => x"ffbf1251",
  1158 => x"70992689",
  1159 => x"38a01270",
  1160 => x"81ff0654",
  1161 => x"51727570",
  1162 => x"81055784",
  1163 => x"808081b7",
  1164 => x"2d811656",
  1165 => x"80748480",
  1166 => x"8080f52d",
  1167 => x"53517171",
  1168 => x"2e833881",
  1169 => x"51758b24",
  1170 => x"853870ff",
  1171 => x"bd388075",
  1172 => x"84808081",
  1173 => x"b72d810b",
  1174 => x"83ffe080",
  1175 => x"0c029805",
  1176 => x"0d0402e0",
  1177 => x"050d797b",
  1178 => x"7d575754",
  1179 => x"80745258",
  1180 => x"8480809f",
  1181 => x"c52d83ff",
  1182 => x"e0800878",
  1183 => x"24527578",
  1184 => x"2e80eb38",
  1185 => x"71782e80",
  1186 => x"e5387478",
  1187 => x"2e80df38",
  1188 => x"83ffe080",
  1189 => x"08148105",
  1190 => x"70848080",
  1191 => x"80f52d54",
  1192 => x"5472782e",
  1193 => x"b938ff15",
  1194 => x"57777725",
  1195 => x"b1387281",
  1196 => x"15ffbf15",
  1197 => x"54555571",
  1198 => x"99268938",
  1199 => x"a0137081",
  1200 => x"ff065652",
  1201 => x"74767081",
  1202 => x"05588480",
  1203 => x"8081b72d",
  1204 => x"81187484",
  1205 => x"808080f5",
  1206 => x"2d545872",
  1207 => x"cc388076",
  1208 => x"84808081",
  1209 => x"b72d8152",
  1210 => x"848080a5",
  1211 => x"f0048052",
  1212 => x"7183ffe0",
  1213 => x"800c02a0",
  1214 => x"050d0402",
  1215 => x"dc050d7a",
  1216 => x"7c7e605b",
  1217 => x"55575280",
  1218 => x"705855af",
  1219 => x"72810509",
  1220 => x"7074079f",
  1221 => x"2a515259",
  1222 => x"75752e81",
  1223 => x"d9388170",
  1224 => x"72065254",
  1225 => x"70752e81",
  1226 => x"cd387281",
  1227 => x"05097074",
  1228 => x"079f2a51",
  1229 => x"51747825",
  1230 => x"81bc3870",
  1231 => x"74065170",
  1232 => x"752e81b2",
  1233 => x"38718480",
  1234 => x"8080f52d",
  1235 => x"5170752e",
  1236 => x"b338fe18",
  1237 => x"54747425",
  1238 => x"ab387081",
  1239 => x"13535770",
  1240 => x"80dc2e09",
  1241 => x"81068338",
  1242 => x"70597673",
  1243 => x"70810555",
  1244 => x"84808081",
  1245 => x"b72d8115",
  1246 => x"72848080",
  1247 => x"80f52d52",
  1248 => x"5570d238",
  1249 => x"7680dc32",
  1250 => x"70810509",
  1251 => x"7072079f",
  1252 => x"2a515252",
  1253 => x"76af2e92",
  1254 => x"3870802e",
  1255 => x"8d387873",
  1256 => x"70810555",
  1257 => x"84808081",
  1258 => x"b72d7584",
  1259 => x"808080f5",
  1260 => x"2d7081ff",
  1261 => x"06525270",
  1262 => x"802eab38",
  1263 => x"ff185474",
  1264 => x"7425a338",
  1265 => x"81165671",
  1266 => x"73708105",
  1267 => x"55848080",
  1268 => x"81b72d81",
  1269 => x"15768480",
  1270 => x"8080f52d",
  1271 => x"7081ff06",
  1272 => x"53535570",
  1273 => x"da388073",
  1274 => x"84808081",
  1275 => x"b72d8151",
  1276 => x"848080a7",
  1277 => x"f8048051",
  1278 => x"7083ffe0",
  1279 => x"800c02a4",
  1280 => x"050d0402",
  1281 => x"fc050d72",
  1282 => x"51807184",
  1283 => x"808081b7",
  1284 => x"2d028405",
  1285 => x"0d0402fc",
  1286 => x"050d728b",
  1287 => x"11848080",
  1288 => x"80f52d70",
  1289 => x"8f06708f",
  1290 => x"32708105",
  1291 => x"09708025",
  1292 => x"83ffe080",
  1293 => x"0c515151",
  1294 => x"51510284",
  1295 => x"050d0402",
  1296 => x"f8050d73",
  1297 => x"8b118480",
  1298 => x"8080f52d",
  1299 => x"5252708f",
  1300 => x"2ea43871",
  1301 => x"84808080",
  1302 => x"f52d5271",
  1303 => x"802e9738",
  1304 => x"7181e52e",
  1305 => x"91387088",
  1306 => x"2e8c3870",
  1307 => x"86065181",
  1308 => x"5270802e",
  1309 => x"83388052",
  1310 => x"7183ffe0",
  1311 => x"800c0288",
  1312 => x"050d0402",
  1313 => x"f8050d73",
  1314 => x"8b118480",
  1315 => x"8080f52d",
  1316 => x"70842a70",
  1317 => x"81065151",
  1318 => x"51518152",
  1319 => x"70833870",
  1320 => x"527183ff",
  1321 => x"e0800c02",
  1322 => x"88050d04",
  1323 => x"02f8050d",
  1324 => x"738b1184",
  1325 => x"808080f5",
  1326 => x"2d70852a",
  1327 => x"70810651",
  1328 => x"51515181",
  1329 => x"52708338",
  1330 => x"70527183",
  1331 => x"ffe0800c",
  1332 => x"0288050d",
  1333 => x"0402fc05",
  1334 => x"0d725180",
  1335 => x"0b84120c",
  1336 => x"80710c02",
  1337 => x"84050d04",
  1338 => x"02f4050d",
  1339 => x"74767008",
  1340 => x"53535370",
  1341 => x"8c388412",
  1342 => x"08730c84",
  1343 => x"8080aa87",
  1344 => x"04841208",
  1345 => x"84120c84",
  1346 => x"12085170",
  1347 => x"8c387108",
  1348 => x"84140c84",
  1349 => x"8080aa9d",
  1350 => x"04710871",
  1351 => x"0c028c05",
  1352 => x"0d0402f0",
  1353 => x"050d7577",
  1354 => x"84120853",
  1355 => x"545470bf",
  1356 => x"38730852",
  1357 => x"71953872",
  1358 => x"740c7284",
  1359 => x"150c7073",
  1360 => x"0c708414",
  1361 => x"0c848080",
  1362 => x"ab900471",
  1363 => x"08730c71",
  1364 => x"84140c71",
  1365 => x"0851708a",
  1366 => x"3872740c",
  1367 => x"848080aa",
  1368 => x"e6047284",
  1369 => x"120c7272",
  1370 => x"0c848080",
  1371 => x"ab900470",
  1372 => x"730c8411",
  1373 => x"0884140c",
  1374 => x"84110852",
  1375 => x"718b3872",
  1376 => x"84150c84",
  1377 => x"8080ab8c",
  1378 => x"0472720c",
  1379 => x"7284120c",
  1380 => x"0290050d",
  1381 => x"0402f405",
  1382 => x"0d88bc15",
  1383 => x"705383ff",
  1384 => x"f2d45253",
  1385 => x"848080a9",
  1386 => x"e82d7252",
  1387 => x"83fff2dc",
  1388 => x"51848080",
  1389 => x"aaa22d02",
  1390 => x"8c050d04",
  1391 => x"02fdb405",
  1392 => x"0d0282d0",
  1393 => x"050883ff",
  1394 => x"e9ec525a",
  1395 => x"848080d1",
  1396 => x"df2d83ff",
  1397 => x"e080087a",
  1398 => x"52568480",
  1399 => x"8099ef2d",
  1400 => x"800b83ff",
  1401 => x"e0800881",
  1402 => x"055a5877",
  1403 => x"792581a0",
  1404 => x"38828454",
  1405 => x"0280c805",
  1406 => x"70547853",
  1407 => x"7a525784",
  1408 => x"80809b9f",
  1409 => x"2d83ffe0",
  1410 => x"8008ff2e",
  1411 => x"09810689",
  1412 => x"38805584",
  1413 => x"8080ad9b",
  1414 => x"0402a805",
  1415 => x"70557754",
  1416 => x"765383ff",
  1417 => x"e9ec5255",
  1418 => x"848080d1",
  1419 => x"f22d83ff",
  1420 => x"e0800880",
  1421 => x"2e903874",
  1422 => x"51848080",
  1423 => x"a9832d83",
  1424 => x"ffe08008",
  1425 => x"8d3883ff",
  1426 => x"e0800855",
  1427 => x"848080ad",
  1428 => x"9b0402bc",
  1429 => x"05848080",
  1430 => x"80e02d70",
  1431 => x"882b83fe",
  1432 => x"80067188",
  1433 => x"2a070288",
  1434 => x"0580c205",
  1435 => x"84808080",
  1436 => x"e02d7088",
  1437 => x"2b83fe80",
  1438 => x"0671882a",
  1439 => x"07728480",
  1440 => x"80290581",
  1441 => x"1c5c5957",
  1442 => x"51578480",
  1443 => x"80abeb04",
  1444 => x"0282d405",
  1445 => x"0876710c",
  1446 => x"55815574",
  1447 => x"83ffe080",
  1448 => x"0c0282cc",
  1449 => x"050d0402",
  1450 => x"ffb8050d",
  1451 => x"83fff2dc",
  1452 => x"08705a56",
  1453 => x"75802e83",
  1454 => x"c8387552",
  1455 => x"83fff2dc",
  1456 => x"51848080",
  1457 => x"a9e82d75",
  1458 => x"5283fff2",
  1459 => x"d4518480",
  1460 => x"80aaa22d",
  1461 => x"f7c41659",
  1462 => x"78802e83",
  1463 => x"a438f7d8",
  1464 => x"165a8284",
  1465 => x"53805279",
  1466 => x"51848080",
  1467 => x"e0f02df9",
  1468 => x"dc165882",
  1469 => x"84538052",
  1470 => x"77518480",
  1471 => x"80e0f02d",
  1472 => x"82845577",
  1473 => x"54828453",
  1474 => x"79526351",
  1475 => x"8480809d",
  1476 => x"ab2d83ff",
  1477 => x"e08008ff",
  1478 => x"2e82ee38",
  1479 => x"83fff2d4",
  1480 => x"08577680",
  1481 => x"2ebd38f7",
  1482 => x"c4175675",
  1483 => x"792eaa38",
  1484 => x"7952f7d8",
  1485 => x"17518480",
  1486 => x"80a0c22d",
  1487 => x"83ffe080",
  1488 => x"08802e95",
  1489 => x"387752f9",
  1490 => x"dc175184",
  1491 => x"8080a0c2",
  1492 => x"2d83ffe0",
  1493 => x"800882b1",
  1494 => x"38841708",
  1495 => x"57848080",
  1496 => x"aea20494",
  1497 => x"19848080",
  1498 => x"80f52d56",
  1499 => x"75993883",
  1500 => x"ffe9ec51",
  1501 => x"848080d1",
  1502 => x"df2d83ff",
  1503 => x"e0800879",
  1504 => x"0c848080",
  1505 => x"afad0478",
  1506 => x"52941951",
  1507 => x"848080ab",
  1508 => x"bc2d83ff",
  1509 => x"e0800856",
  1510 => x"83ffe080",
  1511 => x"088f3878",
  1512 => x"51848080",
  1513 => x"ab952d84",
  1514 => x"8080b193",
  1515 => x"0402a805",
  1516 => x"70558298",
  1517 => x"1a547908",
  1518 => x"5383ffe9",
  1519 => x"ec525684",
  1520 => x"8080d1f2",
  1521 => x"2d83ffe0",
  1522 => x"8008802e",
  1523 => x"81bb3875",
  1524 => x"51848080",
  1525 => x"a9ac2d83",
  1526 => x"ffe08008",
  1527 => x"802e81a9",
  1528 => x"388b5375",
  1529 => x"52849c19",
  1530 => x"51848080",
  1531 => x"ddfd2d61",
  1532 => x"70882b87",
  1533 => x"fc808006",
  1534 => x"7072982b",
  1535 => x"0772882a",
  1536 => x"83fe8006",
  1537 => x"71077398",
  1538 => x"2a078c1d",
  1539 => x"0c515757",
  1540 => x"800b881a",
  1541 => x"0c02bc05",
  1542 => x"84808080",
  1543 => x"e02d7088",
  1544 => x"2b83fe80",
  1545 => x"0671882a",
  1546 => x"07028805",
  1547 => x"80c20584",
  1548 => x"808080e0",
  1549 => x"2d70882b",
  1550 => x"83fe8006",
  1551 => x"71882a07",
  1552 => x"72848080",
  1553 => x"2905841d",
  1554 => x"0c585158",
  1555 => x"ff0b88b0",
  1556 => x"1a0c800b",
  1557 => x"88b41a0c",
  1558 => x"800b901a",
  1559 => x"0cff0b84",
  1560 => x"a81a0cff",
  1561 => x"0b84ac1a",
  1562 => x"0c785283",
  1563 => x"ffe9ec51",
  1564 => x"848080c4",
  1565 => x"9f2d83ff",
  1566 => x"e9ec5184",
  1567 => x"808094a5",
  1568 => x"2d785684",
  1569 => x"8080b193",
  1570 => x"04785184",
  1571 => x"8080ab95",
  1572 => x"2d805675",
  1573 => x"83ffe080",
  1574 => x"0c0280c8",
  1575 => x"050d0402",
  1576 => x"d0050d7d",
  1577 => x"7f6283ff",
  1578 => x"e9ec0b84",
  1579 => x"808080f5",
  1580 => x"2d705672",
  1581 => x"555a5c56",
  1582 => x"59848080",
  1583 => x"e3a82d83",
  1584 => x"ffe08008",
  1585 => x"83ffe080",
  1586 => x"08782976",
  1587 => x"71317c11",
  1588 => x"585d5758",
  1589 => x"76752785",
  1590 => x"38767b31",
  1591 => x"5a84a819",
  1592 => x"08567776",
  1593 => x"2e098106",
  1594 => x"8c3884ac",
  1595 => x"19085684",
  1596 => x"8080b2fd",
  1597 => x"0477802e",
  1598 => x"99388116",
  1599 => x"5577752e",
  1600 => x"0981068e",
  1601 => x"387584ac",
  1602 => x"1a085755",
  1603 => x"848080b2",
  1604 => x"9904800b",
  1605 => x"841a0857",
  1606 => x"55747827",
  1607 => x"80d03802",
  1608 => x"b005fc05",
  1609 => x"54745378",
  1610 => x"5283ffe9",
  1611 => x"ec518480",
  1612 => x"80c4a72d",
  1613 => x"83ffe080",
  1614 => x"08a93875",
  1615 => x"5283ffe9",
  1616 => x"ec518480",
  1617 => x"8094f22d",
  1618 => x"83ffe080",
  1619 => x"085c83ff",
  1620 => x"e0800854",
  1621 => x"74537852",
  1622 => x"83ffe9ec",
  1623 => x"51848080",
  1624 => x"c4af2d7b",
  1625 => x"81165656",
  1626 => x"848080b2",
  1627 => x"990475ff",
  1628 => x"2e933875",
  1629 => x"84ac1a0c",
  1630 => x"7784a81a",
  1631 => x"0c75ff2e",
  1632 => x"09810689",
  1633 => x"38805584",
  1634 => x"8080b3bf",
  1635 => x"04755283",
  1636 => x"ffe9ec51",
  1637 => x"848080cc",
  1638 => x"ca2d7954",
  1639 => x"7f5383ff",
  1640 => x"e080081b",
  1641 => x"5283ffe9",
  1642 => x"ec518480",
  1643 => x"80cda12d",
  1644 => x"795583ff",
  1645 => x"e0800887",
  1646 => x"3883ffe0",
  1647 => x"80085574",
  1648 => x"83ffe080",
  1649 => x"0c02b005",
  1650 => x"0d0402f8",
  1651 => x"050d83ff",
  1652 => x"f2dc5184",
  1653 => x"8080a9d5",
  1654 => x"2d83fff2",
  1655 => x"d4518480",
  1656 => x"80a9d52d",
  1657 => x"83ffe9e4",
  1658 => x"5283fff2",
  1659 => x"dc518480",
  1660 => x"80aaa22d",
  1661 => x"810b83ff",
  1662 => x"e1a00c02",
  1663 => x"88050d04",
  1664 => x"02fc050d",
  1665 => x"83ffeaa8",
  1666 => x"73717084",
  1667 => x"05530c74",
  1668 => x"710c5102",
  1669 => x"84050d04",
  1670 => x"02f4050d",
  1671 => x"83ffe1a0",
  1672 => x"08873884",
  1673 => x"8080b3ca",
  1674 => x"2d7483ff",
  1675 => x"eaa00c75",
  1676 => x"83ffeaa4",
  1677 => x"0c83ffe9",
  1678 => x"ec518480",
  1679 => x"80c4b72d",
  1680 => x"83ffe080",
  1681 => x"085383ff",
  1682 => x"e0800880",
  1683 => x"2e993883",
  1684 => x"ffe08008",
  1685 => x"52848080",
  1686 => x"e8b45184",
  1687 => x"808082e3",
  1688 => x"2d848080",
  1689 => x"b4f40481",
  1690 => x"0b83ffe1",
  1691 => x"a40c83ff",
  1692 => x"e0800853",
  1693 => x"7283ffe0",
  1694 => x"800c028c",
  1695 => x"050d0402",
  1696 => x"f8050d83",
  1697 => x"ffe1a008",
  1698 => x"87388480",
  1699 => x"80b3ca2d",
  1700 => x"83ffeaa8",
  1701 => x"08527180",
  1702 => x"2e833871",
  1703 => x"2d83ffe9",
  1704 => x"ec518480",
  1705 => x"8094a52d",
  1706 => x"83ffeaac",
  1707 => x"08527180",
  1708 => x"2e833871",
  1709 => x"2d028805",
  1710 => x"0d0402e8",
  1711 => x"050d7779",
  1712 => x"56568054",
  1713 => x"83ffe1a0",
  1714 => x"08742e09",
  1715 => x"81068738",
  1716 => x"848080b3",
  1717 => x"ca2d7352",
  1718 => x"83ffe1a4",
  1719 => x"08802e82",
  1720 => x"ff387581",
  1721 => x"05097077",
  1722 => x"07802576",
  1723 => x"81050970",
  1724 => x"78078025",
  1725 => x"72077752",
  1726 => x"52545153",
  1727 => x"7282e138",
  1728 => x"73538480",
  1729 => x"80b7dd04",
  1730 => x"72157084",
  1731 => x"808080f5",
  1732 => x"2d515271",
  1733 => x"80d72e80",
  1734 => x"e8387180",
  1735 => x"d724ad38",
  1736 => x"7180c22e",
  1737 => x"81b03871",
  1738 => x"80c22494",
  1739 => x"3871ab2e",
  1740 => x"80e33871",
  1741 => x"80c12e80",
  1742 => x"d2388480",
  1743 => x"80b7da04",
  1744 => x"7180d22e",
  1745 => x"b2388480",
  1746 => x"80b7da04",
  1747 => x"7180e22e",
  1748 => x"81843871",
  1749 => x"80e2248d",
  1750 => x"387180e1",
  1751 => x"2ead3884",
  1752 => x"8080b7da",
  1753 => x"047180f2",
  1754 => x"2e8d3871",
  1755 => x"80f72e91",
  1756 => x"38848080",
  1757 => x"b7da0473",
  1758 => x"81075484",
  1759 => x"8080b7da",
  1760 => x"0473b207",
  1761 => x"54848080",
  1762 => x"b7da0473",
  1763 => x"a6075484",
  1764 => x"8080b7da",
  1765 => x"04738106",
  1766 => x"5271802e",
  1767 => x"8b387382",
  1768 => x"07548480",
  1769 => x"80b7da04",
  1770 => x"73812a70",
  1771 => x"81065152",
  1772 => x"71802e8b",
  1773 => x"3873b107",
  1774 => x"54848080",
  1775 => x"b7da0473",
  1776 => x"822a7081",
  1777 => x"06515271",
  1778 => x"802e8f38",
  1779 => x"73a70754",
  1780 => x"848080b7",
  1781 => x"da047388",
  1782 => x"07548113",
  1783 => x"53745184",
  1784 => x"8080d8f2",
  1785 => x"2d83ffe0",
  1786 => x"80087324",
  1787 => x"fe9a3880",
  1788 => x"7481d906",
  1789 => x"555383ff",
  1790 => x"eaa40873",
  1791 => x"2e098106",
  1792 => x"86387381",
  1793 => x"d9065483",
  1794 => x"ffeaa808",
  1795 => x"5271802e",
  1796 => x"8338712d",
  1797 => x"73810652",
  1798 => x"719a3873",
  1799 => x"852a7081",
  1800 => x"06515272",
  1801 => x"a2387180",
  1802 => x"2e983873",
  1803 => x"86065271",
  1804 => x"802e8f38",
  1805 => x"75518480",
  1806 => x"80ada72d",
  1807 => x"83ffe080",
  1808 => x"08537280",
  1809 => x"2e8b3873",
  1810 => x"88b81484",
  1811 => x"808081b7",
  1812 => x"2d83ffea",
  1813 => x"ac085271",
  1814 => x"802e8338",
  1815 => x"712d7252",
  1816 => x"7183ffe0",
  1817 => x"800c0298",
  1818 => x"050d0480",
  1819 => x"0b83ffe0",
  1820 => x"800c0402",
  1821 => x"f4050d74",
  1822 => x"5283ffe1",
  1823 => x"a0088738",
  1824 => x"848080b3",
  1825 => x"ca2d7180",
  1826 => x"2e80da38",
  1827 => x"83ffeaa8",
  1828 => x"08537280",
  1829 => x"2e833872",
  1830 => x"2d901208",
  1831 => x"802e8638",
  1832 => x"800b9013",
  1833 => x"0c800b88",
  1834 => x"130c800b",
  1835 => x"8c130c80",
  1836 => x"0b84130c",
  1837 => x"ff0b88b0",
  1838 => x"130c800b",
  1839 => x"88b4130c",
  1840 => x"800b9013",
  1841 => x"0c715184",
  1842 => x"8080ab95",
  1843 => x"2d83ffe9",
  1844 => x"ec518480",
  1845 => x"8094a52d",
  1846 => x"83ffeaac",
  1847 => x"08527180",
  1848 => x"2e833871",
  1849 => x"2d028c05",
  1850 => x"0d0402d0",
  1851 => x"050d7d61",
  1852 => x"6062295a",
  1853 => x"5a5c805b",
  1854 => x"83ffe1a0",
  1855 => x"087b2e09",
  1856 => x"81068738",
  1857 => x"848080b3",
  1858 => x"ca2d7b81",
  1859 => x"0509707d",
  1860 => x"0780257a",
  1861 => x"81050970",
  1862 => x"7c078025",
  1863 => x"72075257",
  1864 => x"5156ff5a",
  1865 => x"7581f238",
  1866 => x"88b81984",
  1867 => x"808080f5",
  1868 => x"2d810655",
  1869 => x"74802e81",
  1870 => x"e0387a5a",
  1871 => x"77802e81",
  1872 => x"d8388819",
  1873 => x"088c1a08",
  1874 => x"5856ff5a",
  1875 => x"75772781",
  1876 => x"c8387716",
  1877 => x"55767527",
  1878 => x"85387676",
  1879 => x"31587589",
  1880 => x"2a7683ff",
  1881 => x"065b5580",
  1882 => x"782581ab",
  1883 => x"387980c4",
  1884 => x"38777b31",
  1885 => x"5683ff76",
  1886 => x"25ba3875",
  1887 => x"80258538",
  1888 => x"83ff1656",
  1889 => x"75892c54",
  1890 => x"7a1c5374",
  1891 => x"52785184",
  1892 => x"8080b19f",
  1893 => x"2d83ffe0",
  1894 => x"8008802e",
  1895 => x"80f93883",
  1896 => x"ffe08008",
  1897 => x"892b83ff",
  1898 => x"e0800816",
  1899 => x"56578480",
  1900 => x"80bc8704",
  1901 => x"88b01908",
  1902 => x"752ea638",
  1903 => x"815484b0",
  1904 => x"19537452",
  1905 => x"78518480",
  1906 => x"80b19f2d",
  1907 => x"83ffe080",
  1908 => x"08802e80",
  1909 => x"c2387488",
  1910 => x"b01a0c80",
  1911 => x"0b88b41a",
  1912 => x"0c84807a",
  1913 => x"31787c31",
  1914 => x"57577577",
  1915 => x"25833875",
  1916 => x"57765379",
  1917 => x"1984b005",
  1918 => x"527a1c51",
  1919 => x"848080dd",
  1920 => x"fd2d8115",
  1921 => x"55805a76",
  1922 => x"1b881a08",
  1923 => x"18881b0c",
  1924 => x"5b777b24",
  1925 => x"fed7387a",
  1926 => x"5a7983ff",
  1927 => x"e0800c02",
  1928 => x"b0050d04",
  1929 => x"02e8050d",
  1930 => x"80029805",
  1931 => x"84808081",
  1932 => x"b72d7754",
  1933 => x"81538152",
  1934 => x"029805fc",
  1935 => x"05518480",
  1936 => x"80b9ea2d",
  1937 => x"83ffe080",
  1938 => x"085583ff",
  1939 => x"e0800881",
  1940 => x"2e098106",
  1941 => x"8b380294",
  1942 => x"05848080",
  1943 => x"80f52d55",
  1944 => x"7483ffe0",
  1945 => x"800c0298",
  1946 => x"050d0402",
  1947 => x"e8050d77",
  1948 => x"797b5853",
  1949 => x"55805372",
  1950 => x"722580d4",
  1951 => x"38ff1254",
  1952 => x"72742580",
  1953 => x"cb387551",
  1954 => x"848080bc",
  1955 => x"a42d800b",
  1956 => x"83ffe080",
  1957 => x"0824a138",
  1958 => x"74135283",
  1959 => x"ffe08008",
  1960 => x"72848080",
  1961 => x"81b72d81",
  1962 => x"135383ff",
  1963 => x"e080088a",
  1964 => x"2e863873",
  1965 => x"7324cf38",
  1966 => x"80732594",
  1967 => x"38721552",
  1968 => x"80728480",
  1969 => x"8081b72d",
  1970 => x"74528480",
  1971 => x"80bdd204",
  1972 => x"80527183",
  1973 => x"ffe0800c",
  1974 => x"0298050d",
  1975 => x"0402e805",
  1976 => x"0d77797b",
  1977 => x"585454ff",
  1978 => x"5583ffe1",
  1979 => x"a0088738",
  1980 => x"848080b3",
  1981 => x"ca2d7452",
  1982 => x"73802e81",
  1983 => x"bc387582",
  1984 => x"32708105",
  1985 => x"09707207",
  1986 => x"80255152",
  1987 => x"5272802e",
  1988 => x"87387452",
  1989 => x"7081a238",
  1990 => x"83ffeaa8",
  1991 => x"08517080",
  1992 => x"2e833870",
  1993 => x"2dff0b88",
  1994 => x"b0150c80",
  1995 => x"0b88b415",
  1996 => x"0c759a38",
  1997 => x"7288150c",
  1998 => x"8c140851",
  1999 => x"70732785",
  2000 => x"38708815",
  2001 => x"0c755584",
  2002 => x"8080bfaa",
  2003 => x"0475812e",
  2004 => x"09810680",
  2005 => x"c5388814",
  2006 => x"08518073",
  2007 => x"249b3872",
  2008 => x"11708816",
  2009 => x"0c8c1508",
  2010 => x"53517171",
  2011 => x"27ba3871",
  2012 => x"88150c84",
  2013 => x"8080bfa8",
  2014 => x"04728105",
  2015 => x"09537073",
  2016 => x"278c3880",
  2017 => x"0b88150c",
  2018 => x"848080bf",
  2019 => x"a8047073",
  2020 => x"3188150c",
  2021 => x"848080bf",
  2022 => x"a8047582",
  2023 => x"2e098106",
  2024 => x"89388c14",
  2025 => x"0888150c",
  2026 => x"805583ff",
  2027 => x"eaac0851",
  2028 => x"70802e83",
  2029 => x"38702d74",
  2030 => x"527183ff",
  2031 => x"e0800c02",
  2032 => x"98050d04",
  2033 => x"02f8050d",
  2034 => x"7352ff51",
  2035 => x"71802ea4",
  2036 => x"3883ffea",
  2037 => x"a8085170",
  2038 => x"802e8338",
  2039 => x"702d7488",
  2040 => x"1308710c",
  2041 => x"5183ffea",
  2042 => x"ac085170",
  2043 => x"802e8338",
  2044 => x"702d8051",
  2045 => x"7083ffe0",
  2046 => x"800c0288",
  2047 => x"050d0402",
  2048 => x"f0050d80",
  2049 => x"54029005",
  2050 => x"fc055275",
  2051 => x"51848080",
  2052 => x"bfc42d73",
  2053 => x"83ffe080",
  2054 => x"0c029005",
  2055 => x"0d0402f8",
  2056 => x"050d7352",
  2057 => x"ff517180",
  2058 => x"2eb13883",
  2059 => x"ffeaa808",
  2060 => x"5170802e",
  2061 => x"8338702d",
  2062 => x"8812088c",
  2063 => x"13083270",
  2064 => x"81050970",
  2065 => x"72079f2a",
  2066 => x"ff1183ff",
  2067 => x"eaac0854",
  2068 => x"51515252",
  2069 => x"71802e83",
  2070 => x"38712d70",
  2071 => x"83ffe080",
  2072 => x"0c028805",
  2073 => x"0d04800b",
  2074 => x"83ffe080",
  2075 => x"0c0402e4",
  2076 => x"050d787a",
  2077 => x"5755ff57",
  2078 => x"83ffe1a0",
  2079 => x"08873884",
  2080 => x"8080b3ca",
  2081 => x"2d83ffea",
  2082 => x"a8085473",
  2083 => x"802e8338",
  2084 => x"732d7451",
  2085 => x"84808099",
  2086 => x"ef2d83ff",
  2087 => x"e08008ff",
  2088 => x"2e098106",
  2089 => x"983883ff",
  2090 => x"e9ec5184",
  2091 => x"8080d1df",
  2092 => x"2d83ffe0",
  2093 => x"80085784",
  2094 => x"8080c1d4",
  2095 => x"04029c05",
  2096 => x"fc055274",
  2097 => x"51848080",
  2098 => x"abbc2d83",
  2099 => x"ffe08008",
  2100 => x"802e9038",
  2101 => x"76537552",
  2102 => x"83ffe9ec",
  2103 => x"51848080",
  2104 => x"d4c12d83",
  2105 => x"ffeaac08",
  2106 => x"5473802e",
  2107 => x"8338732d",
  2108 => x"755476ff",
  2109 => x"2e098106",
  2110 => x"83388054",
  2111 => x"7383ffe0",
  2112 => x"800c029c",
  2113 => x"050d0402",
  2114 => x"ec050d83",
  2115 => x"ffe1a008",
  2116 => x"87388480",
  2117 => x"80b3ca2d",
  2118 => x"83ffeaa8",
  2119 => x"08547380",
  2120 => x"2e833873",
  2121 => x"2d775376",
  2122 => x"5283ffe9",
  2123 => x"ec518480",
  2124 => x"80d4dd2d",
  2125 => x"83ffe080",
  2126 => x"0883ffea",
  2127 => x"ac085555",
  2128 => x"73802e83",
  2129 => x"38732d74",
  2130 => x"83ffe080",
  2131 => x"0c029405",
  2132 => x"0d0402fd",
  2133 => x"cc050d83",
  2134 => x"ffe1a008",
  2135 => x"87388480",
  2136 => x"80b3ca2d",
  2137 => x"83ffeaa8",
  2138 => x"08547380",
  2139 => x"2e833873",
  2140 => x"2d0282a8",
  2141 => x"05705302",
  2142 => x"82bc0508",
  2143 => x"52568480",
  2144 => x"80c0ee2d",
  2145 => x"83ffe080",
  2146 => x"08802e80",
  2147 => x"d5388480",
  2148 => x"80c3cc04",
  2149 => x"02829c05",
  2150 => x"84808080",
  2151 => x"f52d5473",
  2152 => x"802e9538",
  2153 => x"74528480",
  2154 => x"80e8e851",
  2155 => x"84808082",
  2156 => x"e32d8480",
  2157 => x"80c3cc04",
  2158 => x"0282a405",
  2159 => x"08537452",
  2160 => x"848080e8",
  2161 => x"f4518480",
  2162 => x"8082e32d",
  2163 => x"02980570",
  2164 => x"53765255",
  2165 => x"848080c2",
  2166 => x"872d83ff",
  2167 => x"e08008ff",
  2168 => x"b33883ff",
  2169 => x"eaac0854",
  2170 => x"73802e83",
  2171 => x"38732d02",
  2172 => x"82b4050d",
  2173 => x"0402e405",
  2174 => x"0d8002a0",
  2175 => x"05f40553",
  2176 => x"79525384",
  2177 => x"8080c0ee",
  2178 => x"2d83ffe0",
  2179 => x"8008732e",
  2180 => x"83388153",
  2181 => x"7283ffe0",
  2182 => x"800c029c",
  2183 => x"050d0481",
  2184 => x"0b83ffe0",
  2185 => x"800c0480",
  2186 => x"0b83ffe0",
  2187 => x"800c0481",
  2188 => x"0b83ffe0",
  2189 => x"800c0402",
  2190 => x"ffb8050d",
  2191 => x"63578058",
  2192 => x"ff0b84c4",
  2193 => x"180c7784",
  2194 => x"c8180c77",
  2195 => x"a4180c76",
  2196 => x"51848080",
  2197 => x"919d2db4",
  2198 => x"170854ff",
  2199 => x"5573782e",
  2200 => x"87dc3881",
  2201 => x"5380c417",
  2202 => x"70537852",
  2203 => x"59732d83",
  2204 => x"ffe08008",
  2205 => x"782e87c6",
  2206 => x"3884c217",
  2207 => x"84808080",
  2208 => x"e02d54fd",
  2209 => x"557381ab",
  2210 => x"aa2e0981",
  2211 => x"0687af38",
  2212 => x"84c31784",
  2213 => x"808080f5",
  2214 => x"2d84c218",
  2215 => x"84808080",
  2216 => x"f52d7182",
  2217 => x"80290555",
  2218 => x"55fc5573",
  2219 => x"82d4d52e",
  2220 => x"09810687",
  2221 => x"89388486",
  2222 => x"17848080",
  2223 => x"80f52d70",
  2224 => x"81ff0655",
  2225 => x"56738f26",
  2226 => x"a0388174",
  2227 => x"2b7083b0",
  2228 => x"e0065555",
  2229 => x"73782e09",
  2230 => x"81069938",
  2231 => x"74810654",
  2232 => x"73782e09",
  2233 => x"810680d0",
  2234 => x"387581ff",
  2235 => x"06547386",
  2236 => x"2680c538",
  2237 => x"848d1784",
  2238 => x"808080f5",
  2239 => x"2d848c18",
  2240 => x"84808080",
  2241 => x"f52d7181",
  2242 => x"800a2971",
  2243 => x"84808029",
  2244 => x"05848b1a",
  2245 => x"84808080",
  2246 => x"f52d7082",
  2247 => x"80291284",
  2248 => x"8a1c8480",
  2249 => x"8080f52d",
  2250 => x"5574059c",
  2251 => x"1c0c5956",
  2252 => x"56588480",
  2253 => x"80c6bc04",
  2254 => x"779c180c",
  2255 => x"81537852",
  2256 => x"9c170851",
  2257 => x"b4170854",
  2258 => x"732dff55",
  2259 => x"83ffe080",
  2260 => x"08802e85",
  2261 => x"e93880d0",
  2262 => x"17848080",
  2263 => x"80f52d80",
  2264 => x"cf188480",
  2265 => x"8080f52d",
  2266 => x"7072882b",
  2267 => x"0756415f",
  2268 => x"fe557384",
  2269 => x"802e0981",
  2270 => x"0685c338",
  2271 => x"80d11784",
  2272 => x"808080f5",
  2273 => x"2d778480",
  2274 => x"8081b72d",
  2275 => x"80d31784",
  2276 => x"808080f5",
  2277 => x"2d80d218",
  2278 => x"84808080",
  2279 => x"f52d7072",
  2280 => x"882b0780",
  2281 => x"d41a8480",
  2282 => x"8080f52d",
  2283 => x"7081ff06",
  2284 => x"80d61c84",
  2285 => x"808080f5",
  2286 => x"2d80d51d",
  2287 => x"84808080",
  2288 => x"f52d7072",
  2289 => x"882b075b",
  2290 => x"415f5a41",
  2291 => x"5b434173",
  2292 => x"a8188480",
  2293 => x"80818a2d",
  2294 => x"80db1784",
  2295 => x"808080f5",
  2296 => x"2d80da18",
  2297 => x"84808080",
  2298 => x"f52d7072",
  2299 => x"882b0756",
  2300 => x"5e5c7380",
  2301 => x"2e8b3873",
  2302 => x"a0180c84",
  2303 => x"8080c8bf",
  2304 => x"0480eb17",
  2305 => x"84808080",
  2306 => x"f52d80ea",
  2307 => x"18848080",
  2308 => x"80f52d71",
  2309 => x"81800a29",
  2310 => x"71848080",
  2311 => x"290580e9",
  2312 => x"1a848080",
  2313 => x"80f52d70",
  2314 => x"82802912",
  2315 => x"80e81c84",
  2316 => x"808080f5",
  2317 => x"2d547305",
  2318 => x"a01c0c53",
  2319 => x"56595580",
  2320 => x"f3178480",
  2321 => x"8080f52d",
  2322 => x"80f21884",
  2323 => x"808080f5",
  2324 => x"2d718180",
  2325 => x"0a297184",
  2326 => x"80802905",
  2327 => x"80f11a84",
  2328 => x"808080f5",
  2329 => x"2d708280",
  2330 => x"291280f0",
  2331 => x"1c848080",
  2332 => x"80f52d54",
  2333 => x"7305881c",
  2334 => x"0c80f51b",
  2335 => x"84808080",
  2336 => x"f52d80f4",
  2337 => x"1c848080",
  2338 => x"80f52d71",
  2339 => x"82802905",
  2340 => x"53515356",
  2341 => x"59557398",
  2342 => x"18848080",
  2343 => x"818a2d75",
  2344 => x"a0180829",
  2345 => x"701a8c19",
  2346 => x"0ca81884",
  2347 => x"808080e0",
  2348 => x"2d70852b",
  2349 => x"83ff1152",
  2350 => x"58555873",
  2351 => x"80258538",
  2352 => x"87fe1654",
  2353 => x"73892a90",
  2354 => x"180c9c17",
  2355 => x"08197094",
  2356 => x"190c7805",
  2357 => x"84180c84",
  2358 => x"c3178480",
  2359 => x"8080f52d",
  2360 => x"84c21884",
  2361 => x"808080f5",
  2362 => x"2d718280",
  2363 => x"29055555",
  2364 => x"fd557382",
  2365 => x"d4d52e09",
  2366 => x"810682c2",
  2367 => x"3879882b",
  2368 => x"83fe8006",
  2369 => x"7b81ff06",
  2370 => x"7012852b",
  2371 => x"61882b83",
  2372 => x"fe800663",
  2373 => x"81ff0671",
  2374 => x"05705751",
  2375 => x"527105ff",
  2376 => x"05535556",
  2377 => x"848080e2",
  2378 => x"d52d83ff",
  2379 => x"e080087c",
  2380 => x"882b83fe",
  2381 => x"80067e81",
  2382 => x"ff067105",
  2383 => x"705c5155",
  2384 => x"5a73bd38",
  2385 => x"80eb1784",
  2386 => x"808080f5",
  2387 => x"2d80ea18",
  2388 => x"84808080",
  2389 => x"f52d7181",
  2390 => x"800a2971",
  2391 => x"84808029",
  2392 => x"0580e91a",
  2393 => x"84808080",
  2394 => x"f52d7082",
  2395 => x"80291280",
  2396 => x"e81c8480",
  2397 => x"8080f52d",
  2398 => x"5574055d",
  2399 => x"59565658",
  2400 => x"80d81784",
  2401 => x"808080f5",
  2402 => x"2d80d718",
  2403 => x"84808080",
  2404 => x"f52d7182",
  2405 => x"80290570",
  2406 => x"5a555573",
  2407 => x"bd3880e7",
  2408 => x"17848080",
  2409 => x"80f52d80",
  2410 => x"e6188480",
  2411 => x"8080f52d",
  2412 => x"7181800a",
  2413 => x"29718480",
  2414 => x"80290580",
  2415 => x"e51a8480",
  2416 => x"8080f52d",
  2417 => x"70828029",
  2418 => x"1280e41c",
  2419 => x"84808080",
  2420 => x"f52d5473",
  2421 => x"05545956",
  2422 => x"56586088",
  2423 => x"2b83fe80",
  2424 => x"066281ff",
  2425 => x"067f81ff",
  2426 => x"06577105",
  2427 => x"767b2905",
  2428 => x"7971317c",
  2429 => x"31798480",
  2430 => x"8080f52d",
  2431 => x"52585154",
  2432 => x"fb557380",
  2433 => x"2eb83873",
  2434 => x"52755184",
  2435 => x"8080e3a8",
  2436 => x"2d9ff40b",
  2437 => x"83ffe080",
  2438 => x"0827a338",
  2439 => x"83ffe080",
  2440 => x"0883fff4",
  2441 => x"26913880",
  2442 => x"0b88180c",
  2443 => x"800bb018",
  2444 => x"0c848080",
  2445 => x"ccbc0481",
  2446 => x"0bb0180c",
  2447 => x"80557483",
  2448 => x"ffe0800c",
  2449 => x"0280c805",
  2450 => x"0d0402e8",
  2451 => x"050d7779",
  2452 => x"5755b015",
  2453 => x"08af38a8",
  2454 => x"15848080",
  2455 => x"80e02d53",
  2456 => x"72802584",
  2457 => x"388f1353",
  2458 => x"72842a84",
  2459 => x"16080575",
  2460 => x"84808080",
  2461 => x"f52dfe18",
  2462 => x"71297205",
  2463 => x"52565484",
  2464 => x"8080cd96",
  2465 => x"04748480",
  2466 => x"8080f52d",
  2467 => x"fe177129",
  2468 => x"84170805",
  2469 => x"51547383",
  2470 => x"ffe0800c",
  2471 => x"0298050d",
  2472 => x"0402f005",
  2473 => x"0d785377",
  2474 => x"52765175",
  2475 => x"b4110851",
  2476 => x"54732d02",
  2477 => x"90050d04",
  2478 => x"02f0050d",
  2479 => x"78537752",
  2480 => x"765175b8",
  2481 => x"11085154",
  2482 => x"732d0290",
  2483 => x"050d0402",
  2484 => x"d4050d7c",
  2485 => x"7e60625e",
  2486 => x"5c565780",
  2487 => x"705559b0",
  2488 => x"1708792e",
  2489 => x"09810683",
  2490 => x"38815478",
  2491 => x"5874a138",
  2492 => x"73587380",
  2493 => x"2e9a3878",
  2494 => x"55799018",
  2495 => x"082781a0",
  2496 => x"389c1708",
  2497 => x"8c180805",
  2498 => x"1a548480",
  2499 => x"80ceee04",
  2500 => x"74778480",
  2501 => x"8080f52d",
  2502 => x"70547b53",
  2503 => x"55568480",
  2504 => x"80e3a82d",
  2505 => x"83ffe080",
  2506 => x"0874297a",
  2507 => x"71315a54",
  2508 => x"7783ffe0",
  2509 => x"8008279d",
  2510 => x"3883ffe0",
  2511 => x"80085475",
  2512 => x"52765184",
  2513 => x"808094f2",
  2514 => x"2d83ffe0",
  2515 => x"8008ff15",
  2516 => x"555673eb",
  2517 => x"38805575",
  2518 => x"ff2e80c4",
  2519 => x"38755276",
  2520 => x"51848080",
  2521 => x"ccca2d83",
  2522 => x"ffe08008",
  2523 => x"19547a80",
  2524 => x"2e8b3881",
  2525 => x"537a5284",
  2526 => x"8080cf92",
  2527 => x"04815573",
  2528 => x"84c41808",
  2529 => x"2e9a3873",
  2530 => x"84c4180c",
  2531 => x"745380c4",
  2532 => x"17527351",
  2533 => x"b4170854",
  2534 => x"732d83ff",
  2535 => x"e0800855",
  2536 => x"7483ffe0",
  2537 => x"800c02ac",
  2538 => x"050d0402",
  2539 => x"d8050d7b",
  2540 => x"7d7f61b0",
  2541 => x"14087081",
  2542 => x"0509b016",
  2543 => x"08710770",
  2544 => x"09709f2a",
  2545 => x"51515151",
  2546 => x"585c5c59",
  2547 => x"5677bf38",
  2548 => x"81707506",
  2549 => x"55577380",
  2550 => x"2eb43877",
  2551 => x"54799017",
  2552 => x"082780f4",
  2553 => x"389c1608",
  2554 => x"8c170805",
  2555 => x"1ab41708",
  2556 => x"56547880",
  2557 => x"2e8b3876",
  2558 => x"53785284",
  2559 => x"8080d0ce",
  2560 => x"047384c4",
  2561 => x"170c7653",
  2562 => x"848080d0",
  2563 => x"ca04b416",
  2564 => x"08557880",
  2565 => x"2e9c3877",
  2566 => x"52755184",
  2567 => x"8080ccca",
  2568 => x"2d815378",
  2569 => x"5283ffe0",
  2570 => x"80081a51",
  2571 => x"848080d0",
  2572 => x"d0047752",
  2573 => x"75518480",
  2574 => x"80ccca2d",
  2575 => x"83ffe080",
  2576 => x"081a7084",
  2577 => x"c4180c54",
  2578 => x"815380c4",
  2579 => x"16527351",
  2580 => x"742d83ff",
  2581 => x"e0800854",
  2582 => x"7383ffe0",
  2583 => x"800c02a8",
  2584 => x"050d0402",
  2585 => x"f0050d75",
  2586 => x"848080e9",
  2587 => x"84525484",
  2588 => x"808082e3",
  2589 => x"2d848080",
  2590 => x"e99453b0",
  2591 => x"1408812e",
  2592 => x"87388480",
  2593 => x"80e99c53",
  2594 => x"72528480",
  2595 => x"80e9a451",
  2596 => x"84808082",
  2597 => x"e32d8814",
  2598 => x"08528480",
  2599 => x"80e9b051",
  2600 => x"84808082",
  2601 => x"e32d9414",
  2602 => x"08528480",
  2603 => x"80e9d051",
  2604 => x"84808082",
  2605 => x"e32d8414",
  2606 => x"08528480",
  2607 => x"80e9e851",
  2608 => x"84808082",
  2609 => x"e32d7384",
  2610 => x"808080f5",
  2611 => x"2d528480",
  2612 => x"80ea8451",
  2613 => x"84808082",
  2614 => x"e32d0290",
  2615 => x"050d0402",
  2616 => x"fc050d72",
  2617 => x"88110883",
  2618 => x"ffe0800c",
  2619 => x"51028405",
  2620 => x"0d0402ff",
  2621 => x"ac050d66",
  2622 => x"686a4141",
  2623 => x"5e805d81",
  2624 => x"520280d4",
  2625 => x"05ec0551",
  2626 => x"848080a8",
  2627 => x"832d8054",
  2628 => x"7c53811d",
  2629 => x"60537e52",
  2630 => x"5d848080",
  2631 => x"cdcf2d83",
  2632 => x"ffe08008",
  2633 => x"802e828b",
  2634 => x"38805b7a",
  2635 => x"a0291e80",
  2636 => x"c4057052",
  2637 => x"58848080",
  2638 => x"a8bf2d83",
  2639 => x"ffe08008",
  2640 => x"802e81db",
  2641 => x"380280c4",
  2642 => x"05598d53",
  2643 => x"80527851",
  2644 => x"848080e0",
  2645 => x"f02d8057",
  2646 => x"76197719",
  2647 => x"57557584",
  2648 => x"808080f5",
  2649 => x"2d758480",
  2650 => x"8081b72d",
  2651 => x"81177081",
  2652 => x"ff065855",
  2653 => x"877727e0",
  2654 => x"38805a88",
  2655 => x"02840580",
  2656 => x"c5055d57",
  2657 => x"761c7719",
  2658 => x"56567484",
  2659 => x"808080f5",
  2660 => x"2d768480",
  2661 => x"8081b72d",
  2662 => x"74848080",
  2663 => x"80f52d55",
  2664 => x"74a02e83",
  2665 => x"38815a81",
  2666 => x"177081ff",
  2667 => x"0658558a",
  2668 => x"7727d138",
  2669 => x"79802ea2",
  2670 => x"380280c4",
  2671 => x"05848080",
  2672 => x"80f52d55",
  2673 => x"74ae2e92",
  2674 => x"38ae0280",
  2675 => x"d0058480",
  2676 => x"8081b72d",
  2677 => x"848080d3",
  2678 => x"e504a002",
  2679 => x"80d00584",
  2680 => x"808081b7",
  2681 => x"2d7e5278",
  2682 => x"51848080",
  2683 => x"a0c22d83",
  2684 => x"ffe08008",
  2685 => x"802e9538",
  2686 => x"a0537752",
  2687 => x"69518480",
  2688 => x"80ddfd2d",
  2689 => x"81558480",
  2690 => x"80d4b504",
  2691 => x"83ffe080",
  2692 => x"08520280",
  2693 => x"d405ec05",
  2694 => x"51848080",
  2695 => x"a8832d81",
  2696 => x"1b7081ff",
  2697 => x"065c558f",
  2698 => x"7b27fdff",
  2699 => x"38848080",
  2700 => x"d28e0480",
  2701 => x"557483ff",
  2702 => x"e0800c02",
  2703 => x"80d4050d",
  2704 => x"0402fc05",
  2705 => x"0d737584",
  2706 => x"120c5180",
  2707 => x"710c800b",
  2708 => x"88128480",
  2709 => x"8081b72d",
  2710 => x"0284050d",
  2711 => x"0402ffb4",
  2712 => x"050d6466",
  2713 => x"68405b56",
  2714 => x"80520280",
  2715 => x"cc05ec05",
  2716 => x"51848080",
  2717 => x"a8832d80",
  2718 => x"54790853",
  2719 => x"841a0852",
  2720 => x"75518480",
  2721 => x"80cdcf2d",
  2722 => x"83ffe080",
  2723 => x"08802e83",
  2724 => x"d338881a",
  2725 => x"84808080",
  2726 => x"f52d5978",
  2727 => x"8f2683ae",
  2728 => x"3878a029",
  2729 => x"1680c405",
  2730 => x"70525884",
  2731 => x"8080a8bf",
  2732 => x"2d83ffe0",
  2733 => x"8008802e",
  2734 => x"83863880",
  2735 => x"520280cc",
  2736 => x"05ec0551",
  2737 => x"848080a8",
  2738 => x"832d02bc",
  2739 => x"055b8d53",
  2740 => x"80527a51",
  2741 => x"848080e0",
  2742 => x"f02d8057",
  2743 => x"761b7719",
  2744 => x"57557584",
  2745 => x"808080f5",
  2746 => x"2d758480",
  2747 => x"8081b72d",
  2748 => x"81177081",
  2749 => x"ff065855",
  2750 => x"877727e0",
  2751 => x"38805c88",
  2752 => x"028405bd",
  2753 => x"055e5776",
  2754 => x"1d771956",
  2755 => x"56748480",
  2756 => x"8080f52d",
  2757 => x"76848080",
  2758 => x"81b72d74",
  2759 => x"84808080",
  2760 => x"f52d5574",
  2761 => x"a02e8338",
  2762 => x"815c8117",
  2763 => x"7081ff06",
  2764 => x"58558a77",
  2765 => x"27d1387b",
  2766 => x"802ea138",
  2767 => x"02bc0584",
  2768 => x"808080f5",
  2769 => x"2d5574ae",
  2770 => x"2e9238ae",
  2771 => x"0280c805",
  2772 => x"84808081",
  2773 => x"b72d8480",
  2774 => x"80d6e704",
  2775 => x"a00280c8",
  2776 => x"05848080",
  2777 => x"81b72d7a",
  2778 => x"527d5184",
  2779 => x"8080a3fa",
  2780 => x"2d775184",
  2781 => x"8080a983",
  2782 => x"2d83ffe0",
  2783 => x"8008802e",
  2784 => x"9238810b",
  2785 => x"82841f84",
  2786 => x"808081b7",
  2787 => x"2d848080",
  2788 => x"d7a10483",
  2789 => x"ffe08008",
  2790 => x"82841f84",
  2791 => x"808081b7",
  2792 => x"2d9c1884",
  2793 => x"808080f5",
  2794 => x"2d9d1984",
  2795 => x"808080f5",
  2796 => x"2d71982b",
  2797 => x"71902b07",
  2798 => x"9e1b8480",
  2799 => x"8080f52d",
  2800 => x"70882b72",
  2801 => x"079f1d84",
  2802 => x"808080f5",
  2803 => x"2d710770",
  2804 => x"882b87fc",
  2805 => x"80800670",
  2806 => x"72982b07",
  2807 => x"72882a83",
  2808 => x"fe800671",
  2809 => x"0773982a",
  2810 => x"0766828c",
  2811 => x"050c5153",
  2812 => x"51525957",
  2813 => x"951a8480",
  2814 => x"8080f52d",
  2815 => x"941b8480",
  2816 => x"8080f52d",
  2817 => x"71982b71",
  2818 => x"902b079b",
  2819 => x"1d848080",
  2820 => x"80f52d9a",
  2821 => x"1e848080",
  2822 => x"80f52d71",
  2823 => x"882b0772",
  2824 => x"07648288",
  2825 => x"050c811f",
  2826 => x"53555a58",
  2827 => x"515c5774",
  2828 => x"881b8480",
  2829 => x"8081b72d",
  2830 => x"81558480",
  2831 => x"80d8e604",
  2832 => x"81197081",
  2833 => x"ff065a55",
  2834 => x"848080d5",
  2835 => x"9b047908",
  2836 => x"81057a0c",
  2837 => x"800b881b",
  2838 => x"84808081",
  2839 => x"b72d8480",
  2840 => x"80d4f704",
  2841 => x"80557483",
  2842 => x"ffe0800c",
  2843 => x"0280cc05",
  2844 => x"0d0402f4",
  2845 => x"050d7452",
  2846 => x"80727081",
  2847 => x"05548480",
  2848 => x"8080f52d",
  2849 => x"52537073",
  2850 => x"2e933881",
  2851 => x"13727081",
  2852 => x"05548480",
  2853 => x"8080f52d",
  2854 => x"525370ef",
  2855 => x"387283ff",
  2856 => x"e0800c02",
  2857 => x"8c050d04",
  2858 => x"02f0050d",
  2859 => x"75777156",
  2860 => x"54527270",
  2861 => x"81055484",
  2862 => x"808080f5",
  2863 => x"2d517072",
  2864 => x"70810554",
  2865 => x"84808081",
  2866 => x"b72d70e6",
  2867 => x"387383ff",
  2868 => x"e0800c02",
  2869 => x"90050d04",
  2870 => x"02e4050d",
  2871 => x"787a7c72",
  2872 => x"5a545553",
  2873 => x"848080d9",
  2874 => x"f9048114",
  2875 => x"54747370",
  2876 => x"81055584",
  2877 => x"808081b7",
  2878 => x"2d807484",
  2879 => x"808080f5",
  2880 => x"2d7081ff",
  2881 => x"06535656",
  2882 => x"70762e83",
  2883 => x"38815671",
  2884 => x"81050970",
  2885 => x"73079f2a",
  2886 => x"707806ff",
  2887 => x"15555151",
  2888 => x"5170c738",
  2889 => x"71ff2e96",
  2890 => x"38807370",
  2891 => x"81055584",
  2892 => x"808081b7",
  2893 => x"2dff1252",
  2894 => x"848080da",
  2895 => x"a4047683",
  2896 => x"ffe0800c",
  2897 => x"029c050d",
  2898 => x"0402f005",
  2899 => x"0d757771",
  2900 => x"56545271",
  2901 => x"70810553",
  2902 => x"84808080",
  2903 => x"f52d5170",
  2904 => x"f2387270",
  2905 => x"81055484",
  2906 => x"808080f5",
  2907 => x"2d517072",
  2908 => x"70810554",
  2909 => x"84808081",
  2910 => x"b72d70e6",
  2911 => x"387383ff",
  2912 => x"e0800c02",
  2913 => x"90050d04",
  2914 => x"02ec050d",
  2915 => x"76787a72",
  2916 => x"58555552",
  2917 => x"71708105",
  2918 => x"53848080",
  2919 => x"80f52d51",
  2920 => x"70f23884",
  2921 => x"8080dbb7",
  2922 => x"04ff1353",
  2923 => x"72ff2e9a",
  2924 => x"38811281",
  2925 => x"15555273",
  2926 => x"84808080",
  2927 => x"f52d5170",
  2928 => x"72848080",
  2929 => x"81b72d70",
  2930 => x"e0388072",
  2931 => x"84808081",
  2932 => x"b72d7483",
  2933 => x"ffe0800c",
  2934 => x"0294050d",
  2935 => x"0402f005",
  2936 => x"0d757752",
  2937 => x"52848080",
  2938 => x"dc810470",
  2939 => x"84808080",
  2940 => x"f52d5472",
  2941 => x"742e0981",
  2942 => x"06923881",
  2943 => x"12811252",
  2944 => x"52718480",
  2945 => x"8080f52d",
  2946 => x"5372e038",
  2947 => x"71848080",
  2948 => x"80f52d71",
  2949 => x"84808080",
  2950 => x"f52d7171",
  2951 => x"3183ffe0",
  2952 => x"800c5252",
  2953 => x"0290050d",
  2954 => x"0402ec05",
  2955 => x"0d76787a",
  2956 => x"70555354",
  2957 => x"5470802e",
  2958 => x"80c33884",
  2959 => x"8080dccf",
  2960 => x"04ff1151",
  2961 => x"70802ea1",
  2962 => x"38811481",
  2963 => x"14545473",
  2964 => x"84808080",
  2965 => x"f52d5271",
  2966 => x"802e8e38",
  2967 => x"72848080",
  2968 => x"80f52d55",
  2969 => x"71752ed9",
  2970 => x"38738480",
  2971 => x"8080f52d",
  2972 => x"73848080",
  2973 => x"80f52d71",
  2974 => x"71315454",
  2975 => x"547183ff",
  2976 => x"e0800c02",
  2977 => x"94050d04",
  2978 => x"02f4050d",
  2979 => x"74765451",
  2980 => x"848080dd",
  2981 => x"9e047173",
  2982 => x"2e8f3881",
  2983 => x"11517084",
  2984 => x"808080f5",
  2985 => x"2d5271ee",
  2986 => x"387083ff",
  2987 => x"e0800c02",
  2988 => x"8c050d04",
  2989 => x"02ec050d",
  2990 => x"76785653",
  2991 => x"80738480",
  2992 => x"8080f52d",
  2993 => x"7081ff06",
  2994 => x"53535470",
  2995 => x"742ea338",
  2996 => x"7181ff06",
  2997 => x"5170752e",
  2998 => x"09810683",
  2999 => x"38725481",
  3000 => x"13708480",
  3001 => x"8080f52d",
  3002 => x"7081ff06",
  3003 => x"53535370",
  3004 => x"df387383",
  3005 => x"ffe0800c",
  3006 => x"0294050d",
  3007 => x"0402e805",
  3008 => x"0d77797b",
  3009 => x"72720783",
  3010 => x"06545456",
  3011 => x"5670802e",
  3012 => x"aa387476",
  3013 => x"5253ff12",
  3014 => x"5271ff2e",
  3015 => x"80f43872",
  3016 => x"70810554",
  3017 => x"84808080",
  3018 => x"f52d7170",
  3019 => x"81055384",
  3020 => x"808081b7",
  3021 => x"2d848080",
  3022 => x"de960474",
  3023 => x"7673822a",
  3024 => x"ff055354",
  3025 => x"5470ff2e",
  3026 => x"96387370",
  3027 => x"84055508",
  3028 => x"73708405",
  3029 => x"550cff11",
  3030 => x"51848080",
  3031 => x"dec50471",
  3032 => x"fc067016",
  3033 => x"55760572",
  3034 => x"8306ff05",
  3035 => x"525370ff",
  3036 => x"2ea03873",
  3037 => x"70810555",
  3038 => x"84808080",
  3039 => x"f52d7370",
  3040 => x"81055584",
  3041 => x"808081b7",
  3042 => x"2dff1151",
  3043 => x"848080de",
  3044 => x"ee047583",
  3045 => x"ffe0800c",
  3046 => x"0298050d",
  3047 => x"0402f005",
  3048 => x"0d757078",
  3049 => x"ff1b5454",
  3050 => x"545470ff",
  3051 => x"2ea03871",
  3052 => x"70810553",
  3053 => x"84808080",
  3054 => x"f52d7370",
  3055 => x"81055584",
  3056 => x"808081b7",
  3057 => x"2dff1151",
  3058 => x"848080df",
  3059 => x"aa047383",
  3060 => x"ffe0800c",
  3061 => x"0290050d",
  3062 => x"0402ec05",
  3063 => x"0d787779",
  3064 => x"53545284",
  3065 => x"8080dff7",
  3066 => x"04ff1252",
  3067 => x"71ff2e9c",
  3068 => x"38811381",
  3069 => x"12525370",
  3070 => x"84808080",
  3071 => x"f52d7384",
  3072 => x"808080f5",
  3073 => x"2d565473",
  3074 => x"752ede38",
  3075 => x"72848080",
  3076 => x"80f52d71",
  3077 => x"84808080",
  3078 => x"f52d7171",
  3079 => x"3183ffe0",
  3080 => x"800c5253",
  3081 => x"0294050d",
  3082 => x"0402f005",
  3083 => x"0d767877",
  3084 => x"54525384",
  3085 => x"8080e0c4",
  3086 => x"04ff1151",
  3087 => x"70ff2e94",
  3088 => x"38811252",
  3089 => x"71848080",
  3090 => x"80f52d54",
  3091 => x"72742e09",
  3092 => x"8106e638",
  3093 => x"71728480",
  3094 => x"8080f52d",
  3095 => x"53517272",
  3096 => x"2e833880",
  3097 => x"517083ff",
  3098 => x"e0800c02",
  3099 => x"90050d04",
  3100 => x"02f0050d",
  3101 => x"757771ff",
  3102 => x"1b545455",
  3103 => x"5370ff2e",
  3104 => x"96387372",
  3105 => x"70810554",
  3106 => x"84808081",
  3107 => x"b72dff11",
  3108 => x"51848080",
  3109 => x"e0fd0472",
  3110 => x"83ffe080",
  3111 => x"0c029005",
  3112 => x"0d0402f0",
  3113 => x"050d7552",
  3114 => x"848080e1",
  3115 => x"b1048112",
  3116 => x"52807284",
  3117 => x"808080f5",
  3118 => x"2d7081ff",
  3119 => x"06535454",
  3120 => x"70742e83",
  3121 => x"38815470",
  3122 => x"a02e8438",
  3123 => x"73e03872",
  3124 => x"81ff0651",
  3125 => x"70a02e09",
  3126 => x"81069238",
  3127 => x"81127084",
  3128 => x"808080f5",
  3129 => x"2d525284",
  3130 => x"8080e1d4",
  3131 => x"04718480",
  3132 => x"8080f52d",
  3133 => x"70545170",
  3134 => x"802e8338",
  3135 => x"71537283",
  3136 => x"ffe0800c",
  3137 => x"0290050d",
  3138 => x"0402e805",
  3139 => x"0d777957",
  3140 => x"55805473",
  3141 => x"7524b338",
  3142 => x"75742953",
  3143 => x"72752e09",
  3144 => x"81068938",
  3145 => x"80538480",
  3146 => x"80e2ca04",
  3147 => x"74732591",
  3148 => x"38737629",
  3149 => x"76317571",
  3150 => x"31515384",
  3151 => x"8080e2ca",
  3152 => x"04811454",
  3153 => x"848080e2",
  3154 => x"93047283",
  3155 => x"ffe0800c",
  3156 => x"0298050d",
  3157 => x"0402e005",
  3158 => x"0d797b58",
  3159 => x"56807059",
  3160 => x"54775377",
  3161 => x"762eb638",
  3162 => x"77762499",
  3163 => x"38811477",
  3164 => x"19595475",
  3165 => x"7427ea38",
  3166 => x"72547485",
  3167 => x"249f3884",
  3168 => x"8080e39b",
  3169 => x"04737729",
  3170 => x"77317671",
  3171 => x"31902b70",
  3172 => x"902c5156",
  3173 => x"53848080",
  3174 => x"e2f80472",
  3175 => x"547383ff",
  3176 => x"e0800c02",
  3177 => x"a0050d04",
  3178 => x"02f8050d",
  3179 => x"74527351",
  3180 => x"848080e2",
  3181 => x"d52d0288",
  3182 => x"050d0402",
  3183 => x"f8050d74",
  3184 => x"52735184",
  3185 => x"8080e289",
  3186 => x"2d028805",
  3187 => x"0d0402cc",
  3188 => x"050d8480",
  3189 => x"80eaa051",
  3190 => x"84808082",
  3191 => x"e32d8480",
  3192 => x"80eab051",
  3193 => x"84808082",
  3194 => x"e32d8480",
  3195 => x"80eac851",
  3196 => x"84808082",
  3197 => x"e32d8480",
  3198 => x"8087be2d",
  3199 => x"83ffe080",
  3200 => x"08802e95",
  3201 => x"38848080",
  3202 => x"918c2d83",
  3203 => x"ffe08008",
  3204 => x"81065574",
  3205 => x"802e81ce",
  3206 => x"38848080",
  3207 => x"8db72d84",
  3208 => x"8080b3ca",
  3209 => x"2d848080",
  3210 => x"90dc5284",
  3211 => x"808090aa",
  3212 => x"51848080",
  3213 => x"b4982d83",
  3214 => x"ffe08008",
  3215 => x"802e80c4",
  3216 => x"38848080",
  3217 => x"eadc5184",
  3218 => x"808082e3",
  3219 => x"2d815584",
  3220 => x"8080e7b2",
  3221 => x"0483ffe0",
  3222 => x"80085490",
  3223 => x"80805381",
  3224 => x"5280c0c0",
  3225 => x"84518480",
  3226 => x"80b9ea2d",
  3227 => x"83ffe080",
  3228 => x"08528480",
  3229 => x"80eaf851",
  3230 => x"84808082",
  3231 => x"e32d8480",
  3232 => x"80e69504",
  3233 => x"848080eb",
  3234 => x"8c518480",
  3235 => x"8082e32d",
  3236 => x"848080eb",
  3237 => x"a8518480",
  3238 => x"80c2d22d",
  3239 => x"848080eb",
  3240 => x"ac518480",
  3241 => x"8082e32d",
  3242 => x"80538852",
  3243 => x"02a80570",
  3244 => x"52558480",
  3245 => x"8086ae2d",
  3246 => x"848080eb",
  3247 => x"bc527451",
  3248 => x"848080b5",
  3249 => x"ba2d83ff",
  3250 => x"e080085a",
  3251 => x"83ffe080",
  3252 => x"08ff8238",
  3253 => x"848080eb",
  3254 => x"c0518480",
  3255 => x"8082e32d",
  3256 => x"848080e5",
  3257 => x"9c048480",
  3258 => x"80ebdc51",
  3259 => x"84808082",
  3260 => x"e32d7453",
  3261 => x"885202a8",
  3262 => x"05557451",
  3263 => x"84808086",
  3264 => x"ae2d7484",
  3265 => x"8080ec88",
  3266 => x"2e8b3880",
  3267 => x"53885284",
  3268 => x"8080e5fa",
  3269 => x"04805978",
  3270 => x"822b80c0",
  3271 => x"c0871184",
  3272 => x"808080f5",
  3273 => x"2d80c0c0",
  3274 => x"86128480",
  3275 => x"8080f52d",
  3276 => x"71982b71",
  3277 => x"902b0780",
  3278 => x"c0c08514",
  3279 => x"84808080",
  3280 => x"f52d7088",
  3281 => x"2b720780",
  3282 => x"c0c08416",
  3283 => x"84808080",
  3284 => x"f52d7107",
  3285 => x"70882a83",
  3286 => x"fe800670",
  3287 => x"72982a07",
  3288 => x"72882b87",
  3289 => x"fc808006",
  3290 => x"71077398",
  3291 => x"2b07790c",
  3292 => x"51535152",
  3293 => x"53585957",
  3294 => x"58811959",
  3295 => x"83ffff79",
  3296 => x"25ff9438",
  3297 => x"848080ec",
  3298 => x"8c518480",
  3299 => x"8082e32d",
  3300 => x"79518480",
  3301 => x"80b8f32d",
  3302 => x"848080b4",
  3303 => x"ff2d8480",
  3304 => x"8080932d",
  3305 => x"848080ec",
  3306 => x"98518480",
  3307 => x"8082e32d",
  3308 => x"80557483",
  3309 => x"ffe0800c",
  3310 => x"02b4050d",
  3311 => x"04000000",
  3312 => x"00ffffff",
  3313 => x"ff00ffff",
  3314 => x"ffff00ff",
  3315 => x"ffffff00",
  3316 => x"08200800",
  3317 => x"434d4438",
  3318 => x"5f342072",
  3319 => x"6573706f",
  3320 => x"6e73653a",
  3321 => x"2025640a",
  3322 => x"00000000",
  3323 => x"53444843",
  3324 => x"20496e69",
  3325 => x"7469616c",
  3326 => x"697a6174",
  3327 => x"696f6e20",
  3328 => x"6572726f",
  3329 => x"72210a00",
  3330 => x"434d4435",
  3331 => x"38202564",
  3332 => x"0a202000",
  3333 => x"52656164",
  3334 => x"20636f6d",
  3335 => x"6d616e64",
  3336 => x"20666169",
  3337 => x"6c656420",
  3338 => x"61742025",
  3339 => x"64202825",
  3340 => x"64290a00",
  3341 => x"4641545f",
  3342 => x"46533a20",
  3343 => x"4572726f",
  3344 => x"7220636f",
  3345 => x"756c6420",
  3346 => x"6e6f7420",
  3347 => x"6c6f6164",
  3348 => x"20464154",
  3349 => x"20646574",
  3350 => x"61696c73",
  3351 => x"20282564",
  3352 => x"29210d0a",
  3353 => x"00000000",
  3354 => x"2573203c",
  3355 => x"4449523e",
  3356 => x"0d0a0000",
  3357 => x"2573205b",
  3358 => x"25642062",
  3359 => x"79746573",
  3360 => x"5d0d0a00",
  3361 => x"46415420",
  3362 => x"64657461",
  3363 => x"696c733a",
  3364 => x"0d0a0000",
  3365 => x"46415433",
  3366 => x"32000000",
  3367 => x"46415431",
  3368 => x"36000000",
  3369 => x"20547970",
  3370 => x"65203d25",
  3371 => x"73000000",
  3372 => x"20526f6f",
  3373 => x"74204469",
  3374 => x"72204669",
  3375 => x"72737420",
  3376 => x"436c7573",
  3377 => x"74657220",
  3378 => x"3d202578",
  3379 => x"0d0a0000",
  3380 => x"20464154",
  3381 => x"20426567",
  3382 => x"696e204c",
  3383 => x"4241203d",
  3384 => x"20307825",
  3385 => x"780d0a00",
  3386 => x"20436c75",
  3387 => x"73746572",
  3388 => x"20426567",
  3389 => x"696e204c",
  3390 => x"4241203d",
  3391 => x"20307825",
  3392 => x"780d0a00",
  3393 => x"20536563",
  3394 => x"746f7273",
  3395 => x"20506572",
  3396 => x"20436c75",
  3397 => x"73746572",
  3398 => x"203d2025",
  3399 => x"640d0a00",
  3400 => x"426f6f74",
  3401 => x"206f7074",
  3402 => x"696f6e73",
  3403 => x"3a0a0000",
  3404 => x"30203a20",
  3405 => x"426f6f74",
  3406 => x"2066726f",
  3407 => x"6d205344",
  3408 => x"20636172",
  3409 => x"640a0000",
  3410 => x"31203a20",
  3411 => x"426f6f74",
  3412 => x"2066726f",
  3413 => x"6d204a54",
  3414 => x"41470a00",
  3415 => x"4552524f",
  3416 => x"523a204d",
  3417 => x"65646961",
  3418 => x"20617474",
  3419 => x"61636820",
  3420 => x"6661696c",
  3421 => x"65640a00",
  3422 => x"0a202564",
  3423 => x"20627974",
  3424 => x"65732072",
  3425 => x"6561640a",
  3426 => x"00000000",
  3427 => x"4c697374",
  3428 => x"696e6720",
  3429 => x"64697265",
  3430 => x"63746f72",
  3431 => x"6965732e",
  3432 => x"2e2e0a0a",
  3433 => x"00000000",
  3434 => x"2f000000",
  3435 => x"0a415050",
  3436 => x"2046494c",
  3437 => x"45203e3e",
  3438 => x"20000000",
  3439 => x"72620000",
  3440 => x"4552524f",
  3441 => x"523a2052",
  3442 => x"65616420",
  3443 => x"66696c65",
  3444 => x"20666169",
  3445 => x"6c65640a",
  3446 => x"00000000",
  3447 => x"426f6f74",
  3448 => x"696e6720",
  3449 => x"66726f6d",
  3450 => x"204a5441",
  3451 => x"472c2077",
  3452 => x"61697469",
  3453 => x"6e672066",
  3454 => x"6f722075",
  3455 => x"706c6f61",
  3456 => x"6465720a",
  3457 => x"00000000",
  3458 => x"454e4400",
  3459 => x"0a0a456e",
  3460 => x"642e2e2e",
  3461 => x"200a0000",
  3462 => x"73687574",
  3463 => x"646f776e",
  3464 => x"2e0a0000",
others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;

		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end rtl;

