--
-- (C) 2018, ZPUROMGEN, Yosel de Jesus Balibrea Lastre.
--           Automatically Generated ROM file
--           Please do NOT CHANGE!
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity prog_mem is
generic
(
maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
);
port (
		clk : in std_logic;
		areset : in std_logic := '0';
		from_zpu : in ZPU_ToROM;
		to_zpu : out ZPU_FromROM
		);
end prog_mem;

architecture rtl of prog_mem is

	type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

	shared variable ram : ram_type := (
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080e784",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff2",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"8080e3aa",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c32d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870892a",
   171 => x"70810651",
   172 => x"515170f3",
   173 => x"3871c00c",
   174 => x"7183ffe0",
   175 => x"800c0288",
   176 => x"050d0402",
   177 => x"e8050d80",
   178 => x"78575575",
   179 => x"70840557",
   180 => x"08538054",
   181 => x"72982a73",
   182 => x"882b5452",
   183 => x"71802ea0",
   184 => x"38c00870",
   185 => x"892a7081",
   186 => x"06515151",
   187 => x"70f33871",
   188 => x"c00c8115",
   189 => x"81155555",
   190 => x"837425d8",
   191 => x"3871cc38",
   192 => x"7483ffe0",
   193 => x"800c0298",
   194 => x"050d0402",
   195 => x"fc050dc0",
   196 => x"0870882a",
   197 => x"70810651",
   198 => x"515170f3",
   199 => x"38c00870",
   200 => x"81ff0683",
   201 => x"ffe0800c",
   202 => x"51028405",
   203 => x"0d0402e8",
   204 => x"050d777a",
   205 => x"57548055",
   206 => x"84808086",
   207 => x"8b2d83ff",
   208 => x"e0800881",
   209 => x"ff065372",
   210 => x"882e0981",
   211 => x"06a33880",
   212 => x"7525e538",
   213 => x"75802e8d",
   214 => x"38848080",
   215 => x"e7945184",
   216 => x"808085c3",
   217 => x"2dff14ff",
   218 => x"16565484",
   219 => x"808086b8",
   220 => x"04728d2e",
   221 => x"b638e013",
   222 => x"527180de",
   223 => x"26ffb938",
   224 => x"75802e92",
   225 => x"38c00870",
   226 => x"892a7081",
   227 => x"06515152",
   228 => x"71f33872",
   229 => x"c00c7274",
   230 => x"70810556",
   231 => x"84808081",
   232 => x"b72d8115",
   233 => x"55848080",
   234 => x"86b80480",
   235 => x"74848080",
   236 => x"81b72d74",
   237 => x"83ffe080",
   238 => x"0c029805",
   239 => x"0d0402d0",
   240 => x"050d8070",
   241 => x"57578177",
   242 => x"54588852",
   243 => x"02a40570",
   244 => x"52598480",
   245 => x"8086ae2d",
   246 => x"76557419",
   247 => x"70848080",
   248 => x"80f52d89",
   249 => x"0bd01227",
   250 => x"78058118",
   251 => x"58585154",
   252 => x"877525e6",
   253 => x"38807625",
   254 => x"a63802a3",
   255 => x"05557515",
   256 => x"70848080",
   257 => x"80f52dd0",
   258 => x"117a2979",
   259 => x"057a8829",
   260 => x"7b1005ff",
   261 => x"1a5a5b59",
   262 => x"51547580",
   263 => x"24e03876",
   264 => x"83ffe080",
   265 => x"0c02b005",
   266 => x"0d0402f4",
   267 => x"050dd452",
   268 => x"81ff720c",
   269 => x"71085381",
   270 => x"ff720c72",
   271 => x"882b83fe",
   272 => x"80067208",
   273 => x"7081ff06",
   274 => x"51525381",
   275 => x"ff720c72",
   276 => x"7107882b",
   277 => x"72087081",
   278 => x"ff065152",
   279 => x"5381ff72",
   280 => x"0c727107",
   281 => x"882b7208",
   282 => x"7081ff06",
   283 => x"720783ff",
   284 => x"e0800c52",
   285 => x"53028c05",
   286 => x"0d0402f4",
   287 => x"050d7476",
   288 => x"7181ff06",
   289 => x"d40c5353",
   290 => x"83fff2e4",
   291 => x"08853871",
   292 => x"892b5271",
   293 => x"982ad40c",
   294 => x"71902a70",
   295 => x"81ff06d4",
   296 => x"0c517188",
   297 => x"2a7081ff",
   298 => x"06d40c51",
   299 => x"7181ff06",
   300 => x"d40c7290",
   301 => x"2a7081ff",
   302 => x"06d40c51",
   303 => x"d4087081",
   304 => x"ff065151",
   305 => x"82b8bf52",
   306 => x"7081ff2e",
   307 => x"09810694",
   308 => x"3881ff0b",
   309 => x"d40cd408",
   310 => x"7081ff06",
   311 => x"ff145451",
   312 => x"5171e538",
   313 => x"7083ffe0",
   314 => x"800c028c",
   315 => x"050d0402",
   316 => x"fc050d81",
   317 => x"c75181ff",
   318 => x"0bd40cff",
   319 => x"11517080",
   320 => x"25f43802",
   321 => x"84050d04",
   322 => x"02f0050d",
   323 => x"84808089",
   324 => x"ef2d819c",
   325 => x"9f538052",
   326 => x"87fc80f7",
   327 => x"51848080",
   328 => x"88fa2d83",
   329 => x"ffe08008",
   330 => x"5483ffe0",
   331 => x"8008812e",
   332 => x"098106ae",
   333 => x"3881ff0b",
   334 => x"d40c820a",
   335 => x"52849c80",
   336 => x"e9518480",
   337 => x"8088fa2d",
   338 => x"83ffe080",
   339 => x"088e3881",
   340 => x"ff0bd40c",
   341 => x"73538480",
   342 => x"808ae904",
   343 => x"84808089",
   344 => x"ef2dff13",
   345 => x"5372ffae",
   346 => x"387283ff",
   347 => x"e0800c02",
   348 => x"90050d04",
   349 => x"02f4050d",
   350 => x"81ff0bd4",
   351 => x"0c935380",
   352 => x"5287fc80",
   353 => x"c1518480",
   354 => x"8088fa2d",
   355 => x"83ffe080",
   356 => x"088e3881",
   357 => x"ff0bd40c",
   358 => x"81538480",
   359 => x"808bac04",
   360 => x"84808089",
   361 => x"ef2dff13",
   362 => x"5372d438",
   363 => x"7283ffe0",
   364 => x"800c028c",
   365 => x"050d0402",
   366 => x"f0050d84",
   367 => x"808089ef",
   368 => x"2d83aa52",
   369 => x"849c80c8",
   370 => x"51848080",
   371 => x"88fa2d83",
   372 => x"ffe08008",
   373 => x"812e0981",
   374 => x"06a93884",
   375 => x"808088aa",
   376 => x"2d83ffe0",
   377 => x"800883ff",
   378 => x"ff065372",
   379 => x"83aa2ebb",
   380 => x"3883ffe0",
   381 => x"80085284",
   382 => x"8080e798",
   383 => x"51848080",
   384 => x"82e32d84",
   385 => x"80808af4",
   386 => x"2d848080",
   387 => x"8ca30481",
   388 => x"54848080",
   389 => x"8dac0484",
   390 => x"8080e7b0",
   391 => x"51848080",
   392 => x"82e32d80",
   393 => x"54848080",
   394 => x"8dac0481",
   395 => x"ff0bd40c",
   396 => x"b1538480",
   397 => x"808a882d",
   398 => x"83ffe080",
   399 => x"08802e80",
   400 => x"dc388052",
   401 => x"87fc80fa",
   402 => x"51848080",
   403 => x"88fa2d83",
   404 => x"ffe08008",
   405 => x"b63881ff",
   406 => x"0bd40cd4",
   407 => x"085381ff",
   408 => x"0bd40c81",
   409 => x"ff0bd40c",
   410 => x"81ff0bd4",
   411 => x"0c81ff0b",
   412 => x"d40c7286",
   413 => x"2a708106",
   414 => x"83ffe080",
   415 => x"08565153",
   416 => x"72802ea8",
   417 => x"38848080",
   418 => x"8c8f0483",
   419 => x"ffe08008",
   420 => x"52848080",
   421 => x"e7cc5184",
   422 => x"808082e3",
   423 => x"2d72822e",
   424 => x"fef538ff",
   425 => x"135372ff",
   426 => x"89387254",
   427 => x"7383ffe0",
   428 => x"800c0290",
   429 => x"050d0402",
   430 => x"f4050d81",
   431 => x"0b83fff2",
   432 => x"e40cd008",
   433 => x"708f2a70",
   434 => x"81065151",
   435 => x"5372f338",
   436 => x"72d00c84",
   437 => x"808089ef",
   438 => x"2dd00870",
   439 => x"8f2a7081",
   440 => x"06515153",
   441 => x"72f33881",
   442 => x"0bd00c87",
   443 => x"53805284",
   444 => x"d480c051",
   445 => x"84808088",
   446 => x"fa2d83ff",
   447 => x"e0800881",
   448 => x"2e973872",
   449 => x"822e0981",
   450 => x"06893880",
   451 => x"53848080",
   452 => x"8eda04ff",
   453 => x"135372d5",
   454 => x"38848080",
   455 => x"8bb72d83",
   456 => x"ffe08008",
   457 => x"83fff2e4",
   458 => x"0c83ffe0",
   459 => x"80088e38",
   460 => x"815287fc",
   461 => x"80d05184",
   462 => x"808088fa",
   463 => x"2d81ff0b",
   464 => x"d40cd008",
   465 => x"708f2a70",
   466 => x"81065151",
   467 => x"5372f338",
   468 => x"72d00c81",
   469 => x"ff0bd40c",
   470 => x"81537283",
   471 => x"ffe0800c",
   472 => x"028c050d",
   473 => x"04800b83",
   474 => x"ffe0800c",
   475 => x"0402e005",
   476 => x"0d797b57",
   477 => x"57805881",
   478 => x"ff0bd40c",
   479 => x"d008708f",
   480 => x"2a708106",
   481 => x"51515473",
   482 => x"f3388281",
   483 => x"0bd00c81",
   484 => x"ff0bd40c",
   485 => x"765287fc",
   486 => x"80d15184",
   487 => x"808088fa",
   488 => x"2d80dbc6",
   489 => x"df5583ff",
   490 => x"e0800880",
   491 => x"2e9b3883",
   492 => x"ffe08008",
   493 => x"53765284",
   494 => x"8080e7d8",
   495 => x"51848080",
   496 => x"82e32d84",
   497 => x"8080909f",
   498 => x"0481ff0b",
   499 => x"d40cd408",
   500 => x"7081ff06",
   501 => x"51547381",
   502 => x"fe2e0981",
   503 => x"06a53880",
   504 => x"ff548480",
   505 => x"8088aa2d",
   506 => x"83ffe080",
   507 => x"08767084",
   508 => x"05580cff",
   509 => x"14547380",
   510 => x"25e83881",
   511 => x"58848080",
   512 => x"908904ff",
   513 => x"155574c1",
   514 => x"3881ff0b",
   515 => x"d40cd008",
   516 => x"708f2a70",
   517 => x"81065151",
   518 => x"5473f338",
   519 => x"73d00c77",
   520 => x"83ffe080",
   521 => x"0c02a005",
   522 => x"0d0402ec",
   523 => x"050d7678",
   524 => x"7a555555",
   525 => x"80732798",
   526 => x"38735274",
   527 => x"51848080",
   528 => x"8eed2d81",
   529 => x"15848015",
   530 => x"ff155555",
   531 => x"5572ea38",
   532 => x"810b83ff",
   533 => x"e0800c02",
   534 => x"94050d04",
   535 => x"02fc050d",
   536 => x"74518071",
   537 => x"278738ff",
   538 => x"115170fb",
   539 => x"38810b83",
   540 => x"ffe0800c",
   541 => x"0284050d",
   542 => x"0402ec05",
   543 => x"0d765480",
   544 => x"0b84d415",
   545 => x"0cff0b88",
   546 => x"d8150c80",
   547 => x"0b88dc15",
   548 => x"0c84d814",
   549 => x"55848053",
   550 => x"80527451",
   551 => x"848080e0",
   552 => x"cc2d800b",
   553 => x"88e0150c",
   554 => x"84d41408",
   555 => x"88e4150c",
   556 => x"7484d415",
   557 => x"0c029405",
   558 => x"0d0402d8",
   559 => x"050d7b7d",
   560 => x"70565855",
   561 => x"76802e80",
   562 => x"d0388484",
   563 => x"1708802e",
   564 => x"80c538b8",
   565 => x"15085978",
   566 => x"802eb638",
   567 => x"810b8480",
   568 => x"18087094",
   569 => x"18083172",
   570 => x"11a01908",
   571 => x"59575859",
   572 => x"5a747427",
   573 => x"85387476",
   574 => x"315a7953",
   575 => x"76527751",
   576 => x"782d83ff",
   577 => x"e0800854",
   578 => x"83ffe080",
   579 => x"08802e89",
   580 => x"38800b84",
   581 => x"84180c81",
   582 => x"547383ff",
   583 => x"e0800c02",
   584 => x"a8050d04",
   585 => x"02e0050d",
   586 => x"797b5957",
   587 => x"800b84d4",
   588 => x"18085656",
   589 => x"74762e80",
   590 => x"db388480",
   591 => x"15085473",
   592 => x"78268938",
   593 => x"81145473",
   594 => x"7826ae38",
   595 => x"848c1508",
   596 => x"54739638",
   597 => x"75802e8c",
   598 => x"3873848c",
   599 => x"170c8480",
   600 => x"8092e904",
   601 => x"7584d418",
   602 => x"0c74848c",
   603 => x"16085656",
   604 => x"74c83884",
   605 => x"80809394",
   606 => x"0474802e",
   607 => x"97387784",
   608 => x"80160831",
   609 => x"892b7505",
   610 => x"8488160c",
   611 => x"74548480",
   612 => x"8093f604",
   613 => x"84d41708",
   614 => x"848c170c",
   615 => x"7584d418",
   616 => x"0c848416",
   617 => x"08802e9a",
   618 => x"38755276",
   619 => x"51848080",
   620 => x"91ba2d83",
   621 => x"ffe08008",
   622 => x"5483ffe0",
   623 => x"8008802e",
   624 => x"b5387784",
   625 => x"80170c81",
   626 => x"53755284",
   627 => x"80160851",
   628 => x"b4170854",
   629 => x"732d83ff",
   630 => x"e0800893",
   631 => x"38ff0b84",
   632 => x"80170c83",
   633 => x"ffe08008",
   634 => x"54848080",
   635 => x"93f60475",
   636 => x"8488170c",
   637 => x"75547383",
   638 => x"ffe0800c",
   639 => x"02a0050d",
   640 => x"0402f005",
   641 => x"0d7584d4",
   642 => x"11085454",
   643 => x"72802eb1",
   644 => x"38848413",
   645 => x"08802e9e",
   646 => x"38725273",
   647 => x"51848080",
   648 => x"91ba2d83",
   649 => x"ffe08008",
   650 => x"8d3883ff",
   651 => x"e0800853",
   652 => x"84808094",
   653 => x"c304848c",
   654 => x"13085384",
   655 => x"8080948c",
   656 => x"04815372",
   657 => x"83ffe080",
   658 => x"0c029005",
   659 => x"0d0402e8",
   660 => x"050d7779",
   661 => x"55567383",
   662 => x"38825473",
   663 => x"882a53b0",
   664 => x"1608802e",
   665 => x"85387387",
   666 => x"2a539416",
   667 => x"08135275",
   668 => x"51848080",
   669 => x"92a42dff",
   670 => x"5583ffe0",
   671 => x"8008802e",
   672 => x"819a3883",
   673 => x"ffe08008",
   674 => x"84880508",
   675 => x"55b01608",
   676 => x"b2387288",
   677 => x"2b747131",
   678 => x"107083ff",
   679 => x"fe061781",
   680 => x"11848080",
   681 => x"80f52d71",
   682 => x"84808080",
   683 => x"f52d7182",
   684 => x"802905fc",
   685 => x"80881153",
   686 => x"58585151",
   687 => x"53848080",
   688 => x"96930472",
   689 => x"872b7471",
   690 => x"31822b83",
   691 => x"fffc0616",
   692 => x"83118480",
   693 => x"8080f52d",
   694 => x"82128480",
   695 => x"8080f52d",
   696 => x"7181800a",
   697 => x"29718480",
   698 => x"80290581",
   699 => x"14848080",
   700 => x"80f52d70",
   701 => x"82802912",
   702 => x"75848080",
   703 => x"80f52d56",
   704 => x"7505f00a",
   705 => x"06ff8080",
   706 => x"80881153",
   707 => x"55535459",
   708 => x"575553ff",
   709 => x"55877327",
   710 => x"83387355",
   711 => x"7483ffe0",
   712 => x"800c0298",
   713 => x"050d0402",
   714 => x"e0050d79",
   715 => x"7b5856b0",
   716 => x"1608802e",
   717 => x"81ba3898",
   718 => x"16848080",
   719 => x"80e02d9c",
   720 => x"17080552",
   721 => x"75518480",
   722 => x"8092a42d",
   723 => x"83ffe080",
   724 => x"085883ff",
   725 => x"e0800880",
   726 => x"2e819538",
   727 => x"83ffe080",
   728 => x"08848805",
   729 => x"08547683",
   730 => x"ec158480",
   731 => x"8081b72d",
   732 => x"83ffe080",
   733 => x"08848805",
   734 => x"0877882a",
   735 => x"55557383",
   736 => x"ed168480",
   737 => x"8081b72d",
   738 => x"83ffe080",
   739 => x"08848805",
   740 => x"0877902a",
   741 => x"55557383",
   742 => x"ee168480",
   743 => x"8081b72d",
   744 => x"83ffe080",
   745 => x"08848805",
   746 => x"0877982a",
   747 => x"55557383",
   748 => x"ef168480",
   749 => x"8081b72d",
   750 => x"810b83ff",
   751 => x"e0800884",
   752 => x"84050c76",
   753 => x"a4170cb8",
   754 => x"16085473",
   755 => x"802e9538",
   756 => x"815383ff",
   757 => x"e0800852",
   758 => x"83ffe080",
   759 => x"08848005",
   760 => x"0851732d",
   761 => x"ff0b8480",
   762 => x"190c800b",
   763 => x"8484190c",
   764 => x"02a0050d",
   765 => x"0402d005",
   766 => x"0d7d5780",
   767 => x"705956a0",
   768 => x"1708762e",
   769 => x"81ba3894",
   770 => x"17081852",
   771 => x"76518480",
   772 => x"8092a42d",
   773 => x"83ffe080",
   774 => x"08802e81",
   775 => x"a338800b",
   776 => x"b0180883",
   777 => x"ffe08008",
   778 => x"84880508",
   779 => x"5b5b5574",
   780 => x"83ffff06",
   781 => x"5379ad38",
   782 => x"72198111",
   783 => x"84808080",
   784 => x"f52d7184",
   785 => x"808080f5",
   786 => x"2d718280",
   787 => x"29057081",
   788 => x"05097080",
   789 => x"251a821a",
   790 => x"5a5a5152",
   791 => x"55538480",
   792 => x"8099ae04",
   793 => x"72198311",
   794 => x"84808080",
   795 => x"f52d8212",
   796 => x"84808080",
   797 => x"f52d7181",
   798 => x"800a2971",
   799 => x"84808029",
   800 => x"05811484",
   801 => x"808080f5",
   802 => x"2d708280",
   803 => x"29127584",
   804 => x"808080f5",
   805 => x"2d710570",
   806 => x"81050970",
   807 => x"72078025",
   808 => x"7e05841e",
   809 => x"5e5e5751",
   810 => x"5253575d",
   811 => x"5d5383ff",
   812 => x"7527fefb",
   813 => x"38811858",
   814 => x"a0170878",
   815 => x"26fec838",
   816 => x"7583ffe0",
   817 => x"800c02b0",
   818 => x"050d0402",
   819 => x"ec050d76",
   820 => x"538054ff",
   821 => x"5272742e",
   822 => x"81963872",
   823 => x"84808080",
   824 => x"f52d5170",
   825 => x"af2e0981",
   826 => x"068c3870",
   827 => x"81145455",
   828 => x"8480809a",
   829 => x"a0048113",
   830 => x"84808080",
   831 => x"f52d5170",
   832 => x"ba2e9638",
   833 => x"82138480",
   834 => x"8080f52d",
   835 => x"51ff5270",
   836 => x"80dc2e09",
   837 => x"810680d8",
   838 => x"3880dc0b",
   839 => x"83145455",
   840 => x"72848080",
   841 => x"80f52d70",
   842 => x"81ff0652",
   843 => x"5270802e",
   844 => x"bc387181",
   845 => x"ff065170",
   846 => x"802ea938",
   847 => x"7181ff06",
   848 => x"81145351",
   849 => x"70752e09",
   850 => x"81068938",
   851 => x"71538480",
   852 => x"809ae404",
   853 => x"71728480",
   854 => x"8080f52d",
   855 => x"53538480",
   856 => x"809ab204",
   857 => x"81145484",
   858 => x"80809aa0",
   859 => x"04ff1452",
   860 => x"7183ffe0",
   861 => x"800c0294",
   862 => x"050d0402",
   863 => x"d0050d7d",
   864 => x"7f616358",
   865 => x"5d5d5380",
   866 => x"70748105",
   867 => x"09707607",
   868 => x"73257074",
   869 => x"7a250751",
   870 => x"51545b58",
   871 => x"ff547178",
   872 => x"2e098106",
   873 => x"81d63872",
   874 => x"84808080",
   875 => x"f52d5271",
   876 => x"af2e0981",
   877 => x"068c3871",
   878 => x"81145457",
   879 => x"8480809b",
   880 => x"ec048113",
   881 => x"84808080",
   882 => x"f52d5271",
   883 => x"ba2e9638",
   884 => x"82138480",
   885 => x"8080f52d",
   886 => x"52ff5471",
   887 => x"80dc2e09",
   888 => x"81068198",
   889 => x"3880dc0b",
   890 => x"83145457",
   891 => x"72518480",
   892 => x"80d8ce2d",
   893 => x"800b83ff",
   894 => x"e0800825",
   895 => x"80cf38ff",
   896 => x"1583ffe0",
   897 => x"80085559",
   898 => x"72848080",
   899 => x"80f52d70",
   900 => x"81ff0670",
   901 => x"79327081",
   902 => x"05097080",
   903 => x"251e5e51",
   904 => x"54565679",
   905 => x"7c2e0981",
   906 => x"06993874",
   907 => x"772e9438",
   908 => x"7779258f",
   909 => x"387a1852",
   910 => x"75728480",
   911 => x"8081b72d",
   912 => x"81185881",
   913 => x"13ff1555",
   914 => x"5373ffbc",
   915 => x"387a8480",
   916 => x"8080f52d",
   917 => x"5271802e",
   918 => x"95388480",
   919 => x"80eae851",
   920 => x"84808085",
   921 => x"c32d8054",
   922 => x"8480809c",
   923 => x"fc048480",
   924 => x"80eae851",
   925 => x"84808085",
   926 => x"c32dff54",
   927 => x"7383ffe0",
   928 => x"800c02b0",
   929 => x"050d0402",
   930 => x"d8050d7b",
   931 => x"7d7f6173",
   932 => x"555c5c59",
   933 => x"57848080",
   934 => x"99cb2d83",
   935 => x"ffe08008",
   936 => x"83ffe080",
   937 => x"08565683",
   938 => x"ffe08008",
   939 => x"ff2e80f2",
   940 => x"387f5478",
   941 => x"5383ffe0",
   942 => x"80085276",
   943 => x"51848080",
   944 => x"9afb2dff",
   945 => x"5583ffe0",
   946 => x"800880d6",
   947 => x"38759338",
   948 => x"83ffe080",
   949 => x"08788480",
   950 => x"8081b72d",
   951 => x"8480809e",
   952 => x"a0047651",
   953 => x"848080d8",
   954 => x"ce2d83ff",
   955 => x"e0800879",
   956 => x"52558480",
   957 => x"80d8ce2d",
   958 => x"7483ffe0",
   959 => x"80083155",
   960 => x"79752583",
   961 => x"38795574",
   962 => x"53765277",
   963 => x"51848080",
   964 => x"ddd92d74",
   965 => x"18ff0555",
   966 => x"80758480",
   967 => x"8081b72d",
   968 => x"80557483",
   969 => x"ffe0800c",
   970 => x"02a8050d",
   971 => x"0402e005",
   972 => x"0d797bff",
   973 => x"1e565657",
   974 => x"73ff2e80",
   975 => x"d7387684",
   976 => x"808080f5",
   977 => x"2d707684",
   978 => x"808080f5",
   979 => x"2d70ffbf",
   980 => x"14555954",
   981 => x"59537099",
   982 => x"268938a0",
   983 => x"137081ff",
   984 => x"065951ff",
   985 => x"bf125170",
   986 => x"99268938",
   987 => x"a0127081",
   988 => x"ff065751",
   989 => x"77763151",
   990 => x"709c3872",
   991 => x"802e9538",
   992 => x"71802e90",
   993 => x"38811781",
   994 => x"16ff1656",
   995 => x"56578480",
   996 => x"809eb804",
   997 => x"80517083",
   998 => x"ffe0800c",
   999 => x"02a0050d",
  1000 => x"0402ec05",
  1001 => x"0d7654ff",
  1002 => x"74545572",
  1003 => x"84808080",
  1004 => x"f52d7081",
  1005 => x"ff065252",
  1006 => x"70802e9b",
  1007 => x"387181ff",
  1008 => x"065170ae",
  1009 => x"2e098106",
  1010 => x"85387274",
  1011 => x"31558113",
  1012 => x"53848080",
  1013 => x"9fab0474",
  1014 => x"83ffe080",
  1015 => x"0c029405",
  1016 => x"0d0402ec",
  1017 => x"050d7678",
  1018 => x"707113ff",
  1019 => x"05555555",
  1020 => x"5573802e",
  1021 => x"9e387184",
  1022 => x"808080f5",
  1023 => x"2d5170a0",
  1024 => x"2e098106",
  1025 => x"8e387175",
  1026 => x"31ff13ff",
  1027 => x"16565353",
  1028 => x"73e43872",
  1029 => x"83ffe080",
  1030 => x"0c029405",
  1031 => x"0d0402d4",
  1032 => x"050d7c7e",
  1033 => x"59598079",
  1034 => x"52578480",
  1035 => x"809fa12d",
  1036 => x"83ffe080",
  1037 => x"08785256",
  1038 => x"8480809f",
  1039 => x"a12d83ff",
  1040 => x"e0800876",
  1041 => x"09708105",
  1042 => x"09707207",
  1043 => x"7a255156",
  1044 => x"565a83ff",
  1045 => x"e08008ff",
  1046 => x"2e8c3876",
  1047 => x"5b73772e",
  1048 => x"09810681",
  1049 => x"f73883ff",
  1050 => x"e0800809",
  1051 => x"70810509",
  1052 => x"70720780",
  1053 => x"25515555",
  1054 => x"75ff2e80",
  1055 => x"e238805b",
  1056 => x"737b2e09",
  1057 => x"810681d4",
  1058 => x"3875ff2e",
  1059 => x"80d13875",
  1060 => x"19810583",
  1061 => x"ffe08008",
  1062 => x"19810571",
  1063 => x"53565784",
  1064 => x"8080d8ce",
  1065 => x"2d83ffe0",
  1066 => x"80087552",
  1067 => x"54848080",
  1068 => x"d8ce2d73",
  1069 => x"83ffe080",
  1070 => x"082e0981",
  1071 => x"06819d38",
  1072 => x"73537452",
  1073 => x"76518480",
  1074 => x"809ead2d",
  1075 => x"757a5555",
  1076 => x"83ffe080",
  1077 => x"087b2ea3",
  1078 => x"38848080",
  1079 => x"a2dc0478",
  1080 => x"51848080",
  1081 => x"d8ce2d83",
  1082 => x"ffe08008",
  1083 => x"78525584",
  1084 => x"8080d8ce",
  1085 => x"2d83ffe0",
  1086 => x"80085474",
  1087 => x"52785184",
  1088 => x"80809fe2",
  1089 => x"2d83ffe0",
  1090 => x"80087453",
  1091 => x"78525584",
  1092 => x"80809fe2",
  1093 => x"2d805b74",
  1094 => x"83ffe080",
  1095 => x"082e0981",
  1096 => x"06ba3883",
  1097 => x"ffe08008",
  1098 => x"53775278",
  1099 => x"51848080",
  1100 => x"9ead2d83",
  1101 => x"ffe08008",
  1102 => x"7b2e9338",
  1103 => x"848080ea",
  1104 => x"e8518480",
  1105 => x"8085c32d",
  1106 => x"848080a2",
  1107 => x"dc048480",
  1108 => x"80eae851",
  1109 => x"84808085",
  1110 => x"c32d815b",
  1111 => x"7a83ffe0",
  1112 => x"800c02ac",
  1113 => x"050d0402",
  1114 => x"f0050d75",
  1115 => x"5372802e",
  1116 => x"80d73872",
  1117 => x"84808080",
  1118 => x"f52d7081",
  1119 => x"ff065252",
  1120 => x"70802e80",
  1121 => x"c4388113",
  1122 => x"84808080",
  1123 => x"f52d5170",
  1124 => x"af387072",
  1125 => x"81ff0652",
  1126 => x"547080dc",
  1127 => x"2e098106",
  1128 => x"83388154",
  1129 => x"70af3270",
  1130 => x"81050970",
  1131 => x"80257607",
  1132 => x"51515170",
  1133 => x"802e8938",
  1134 => x"81518480",
  1135 => x"80a3cb04",
  1136 => x"81135384",
  1137 => x"8080a2f3",
  1138 => x"04805170",
  1139 => x"83ffe080",
  1140 => x"0c029005",
  1141 => x"0d0402e8",
  1142 => x"050d7779",
  1143 => x"55558056",
  1144 => x"848080a4",
  1145 => x"90047181",
  1146 => x"15555371",
  1147 => x"a02ea138",
  1148 => x"ffbf1251",
  1149 => x"70992689",
  1150 => x"38a01270",
  1151 => x"81ff0654",
  1152 => x"51727570",
  1153 => x"81055784",
  1154 => x"808081b7",
  1155 => x"2d811656",
  1156 => x"80748480",
  1157 => x"8080f52d",
  1158 => x"53517171",
  1159 => x"2e833881",
  1160 => x"51758b24",
  1161 => x"853870ff",
  1162 => x"bd388075",
  1163 => x"84808081",
  1164 => x"b72d810b",
  1165 => x"83ffe080",
  1166 => x"0c029805",
  1167 => x"0d0402e0",
  1168 => x"050d797b",
  1169 => x"7d575754",
  1170 => x"80745258",
  1171 => x"8480809f",
  1172 => x"a12d83ff",
  1173 => x"e0800878",
  1174 => x"24527578",
  1175 => x"2e80eb38",
  1176 => x"71782e80",
  1177 => x"e5387478",
  1178 => x"2e80df38",
  1179 => x"83ffe080",
  1180 => x"08148105",
  1181 => x"70848080",
  1182 => x"80f52d54",
  1183 => x"5472782e",
  1184 => x"b938ff15",
  1185 => x"57777725",
  1186 => x"b1387281",
  1187 => x"15ffbf15",
  1188 => x"54555571",
  1189 => x"99268938",
  1190 => x"a0137081",
  1191 => x"ff065652",
  1192 => x"74767081",
  1193 => x"05588480",
  1194 => x"8081b72d",
  1195 => x"81187484",
  1196 => x"808080f5",
  1197 => x"2d545872",
  1198 => x"cc388076",
  1199 => x"84808081",
  1200 => x"b72d8152",
  1201 => x"848080a5",
  1202 => x"cc048052",
  1203 => x"7183ffe0",
  1204 => x"800c02a0",
  1205 => x"050d0402",
  1206 => x"dc050d7a",
  1207 => x"7c7e605b",
  1208 => x"55575280",
  1209 => x"705855af",
  1210 => x"72810509",
  1211 => x"7074079f",
  1212 => x"2a515259",
  1213 => x"75752e81",
  1214 => x"d9388170",
  1215 => x"72065254",
  1216 => x"70752e81",
  1217 => x"cd387281",
  1218 => x"05097074",
  1219 => x"079f2a51",
  1220 => x"51747825",
  1221 => x"81bc3870",
  1222 => x"74065170",
  1223 => x"752e81b2",
  1224 => x"38718480",
  1225 => x"8080f52d",
  1226 => x"5170752e",
  1227 => x"b338fe18",
  1228 => x"54747425",
  1229 => x"ab387081",
  1230 => x"13535770",
  1231 => x"80dc2e09",
  1232 => x"81068338",
  1233 => x"70597673",
  1234 => x"70810555",
  1235 => x"84808081",
  1236 => x"b72d8115",
  1237 => x"72848080",
  1238 => x"80f52d52",
  1239 => x"5570d238",
  1240 => x"7680dc32",
  1241 => x"70810509",
  1242 => x"7072079f",
  1243 => x"2a515252",
  1244 => x"76af2e92",
  1245 => x"3870802e",
  1246 => x"8d387873",
  1247 => x"70810555",
  1248 => x"84808081",
  1249 => x"b72d7584",
  1250 => x"808080f5",
  1251 => x"2d7081ff",
  1252 => x"06525270",
  1253 => x"802eab38",
  1254 => x"ff185474",
  1255 => x"7425a338",
  1256 => x"81165671",
  1257 => x"73708105",
  1258 => x"55848080",
  1259 => x"81b72d81",
  1260 => x"15768480",
  1261 => x"8080f52d",
  1262 => x"7081ff06",
  1263 => x"53535570",
  1264 => x"da388073",
  1265 => x"84808081",
  1266 => x"b72d8151",
  1267 => x"848080a7",
  1268 => x"d4048051",
  1269 => x"7083ffe0",
  1270 => x"800c02a4",
  1271 => x"050d0402",
  1272 => x"fc050d72",
  1273 => x"51807184",
  1274 => x"808081b7",
  1275 => x"2d028405",
  1276 => x"0d0402fc",
  1277 => x"050d728b",
  1278 => x"11848080",
  1279 => x"80f52d70",
  1280 => x"8f06708f",
  1281 => x"32708105",
  1282 => x"09708025",
  1283 => x"83ffe080",
  1284 => x"0c515151",
  1285 => x"51510284",
  1286 => x"050d0402",
  1287 => x"f8050d73",
  1288 => x"8b118480",
  1289 => x"8080f52d",
  1290 => x"5252708f",
  1291 => x"2ea43871",
  1292 => x"84808080",
  1293 => x"f52d5271",
  1294 => x"802e9738",
  1295 => x"7181e52e",
  1296 => x"91387088",
  1297 => x"2e8c3870",
  1298 => x"86065181",
  1299 => x"5270802e",
  1300 => x"83388052",
  1301 => x"7183ffe0",
  1302 => x"800c0288",
  1303 => x"050d0402",
  1304 => x"f8050d73",
  1305 => x"8b118480",
  1306 => x"8080f52d",
  1307 => x"70842a70",
  1308 => x"81065151",
  1309 => x"51518152",
  1310 => x"70833870",
  1311 => x"527183ff",
  1312 => x"e0800c02",
  1313 => x"88050d04",
  1314 => x"02f8050d",
  1315 => x"738b1184",
  1316 => x"808080f5",
  1317 => x"2d70852a",
  1318 => x"70810651",
  1319 => x"51515181",
  1320 => x"52708338",
  1321 => x"70527183",
  1322 => x"ffe0800c",
  1323 => x"0288050d",
  1324 => x"0402fc05",
  1325 => x"0d725180",
  1326 => x"0b84120c",
  1327 => x"80710c02",
  1328 => x"84050d04",
  1329 => x"02f4050d",
  1330 => x"74767008",
  1331 => x"53535370",
  1332 => x"8c388412",
  1333 => x"08730c84",
  1334 => x"8080a9e3",
  1335 => x"04841208",
  1336 => x"84120c84",
  1337 => x"12085170",
  1338 => x"8c387108",
  1339 => x"84140c84",
  1340 => x"8080a9f9",
  1341 => x"04710871",
  1342 => x"0c028c05",
  1343 => x"0d0402f0",
  1344 => x"050d7577",
  1345 => x"84120853",
  1346 => x"545470bf",
  1347 => x"38730852",
  1348 => x"71953872",
  1349 => x"740c7284",
  1350 => x"150c7073",
  1351 => x"0c708414",
  1352 => x"0c848080",
  1353 => x"aaec0471",
  1354 => x"08730c71",
  1355 => x"84140c71",
  1356 => x"0851708a",
  1357 => x"3872740c",
  1358 => x"848080aa",
  1359 => x"c2047284",
  1360 => x"120c7272",
  1361 => x"0c848080",
  1362 => x"aaec0470",
  1363 => x"730c8411",
  1364 => x"0884140c",
  1365 => x"84110852",
  1366 => x"718b3872",
  1367 => x"84150c84",
  1368 => x"8080aae8",
  1369 => x"0472720c",
  1370 => x"7284120c",
  1371 => x"0290050d",
  1372 => x"0402f405",
  1373 => x"0d88bc15",
  1374 => x"705383ff",
  1375 => x"f2d45253",
  1376 => x"848080a9",
  1377 => x"c42d7252",
  1378 => x"83fff2dc",
  1379 => x"51848080",
  1380 => x"a9fe2d02",
  1381 => x"8c050d04",
  1382 => x"02fdb405",
  1383 => x"0d0282d0",
  1384 => x"050883ff",
  1385 => x"e9ec525a",
  1386 => x"848080d1",
  1387 => x"bb2d83ff",
  1388 => x"e080087a",
  1389 => x"52568480",
  1390 => x"8099cb2d",
  1391 => x"800b83ff",
  1392 => x"e0800881",
  1393 => x"055a5877",
  1394 => x"792581a0",
  1395 => x"38828454",
  1396 => x"0280c805",
  1397 => x"70547853",
  1398 => x"7a525784",
  1399 => x"80809afb",
  1400 => x"2d83ffe0",
  1401 => x"8008ff2e",
  1402 => x"09810689",
  1403 => x"38805584",
  1404 => x"8080acf7",
  1405 => x"0402a805",
  1406 => x"70557754",
  1407 => x"765383ff",
  1408 => x"e9ec5255",
  1409 => x"848080d1",
  1410 => x"ce2d83ff",
  1411 => x"e0800880",
  1412 => x"2e903874",
  1413 => x"51848080",
  1414 => x"a8df2d83",
  1415 => x"ffe08008",
  1416 => x"8d3883ff",
  1417 => x"e0800855",
  1418 => x"848080ac",
  1419 => x"f70402bc",
  1420 => x"05848080",
  1421 => x"80e02d70",
  1422 => x"882b83fe",
  1423 => x"80067188",
  1424 => x"2a070288",
  1425 => x"0580c205",
  1426 => x"84808080",
  1427 => x"e02d7088",
  1428 => x"2b83fe80",
  1429 => x"0671882a",
  1430 => x"07728480",
  1431 => x"80290581",
  1432 => x"1c5c5957",
  1433 => x"51578480",
  1434 => x"80abc704",
  1435 => x"0282d405",
  1436 => x"0876710c",
  1437 => x"55815574",
  1438 => x"83ffe080",
  1439 => x"0c0282cc",
  1440 => x"050d0402",
  1441 => x"ffb8050d",
  1442 => x"83fff2dc",
  1443 => x"08705a56",
  1444 => x"75802e83",
  1445 => x"c8387552",
  1446 => x"83fff2dc",
  1447 => x"51848080",
  1448 => x"a9c42d75",
  1449 => x"5283fff2",
  1450 => x"d4518480",
  1451 => x"80a9fe2d",
  1452 => x"f7c41659",
  1453 => x"78802e83",
  1454 => x"a438f7d8",
  1455 => x"165a8284",
  1456 => x"53805279",
  1457 => x"51848080",
  1458 => x"e0cc2df9",
  1459 => x"dc165882",
  1460 => x"84538052",
  1461 => x"77518480",
  1462 => x"80e0cc2d",
  1463 => x"82845577",
  1464 => x"54828453",
  1465 => x"79526351",
  1466 => x"8480809d",
  1467 => x"872d83ff",
  1468 => x"e08008ff",
  1469 => x"2e82ee38",
  1470 => x"83fff2d4",
  1471 => x"08577680",
  1472 => x"2ebd38f7",
  1473 => x"c4175675",
  1474 => x"792eaa38",
  1475 => x"7952f7d8",
  1476 => x"17518480",
  1477 => x"80a09e2d",
  1478 => x"83ffe080",
  1479 => x"08802e95",
  1480 => x"387752f9",
  1481 => x"dc175184",
  1482 => x"8080a09e",
  1483 => x"2d83ffe0",
  1484 => x"800882b1",
  1485 => x"38841708",
  1486 => x"57848080",
  1487 => x"adfe0494",
  1488 => x"19848080",
  1489 => x"80f52d56",
  1490 => x"75993883",
  1491 => x"ffe9ec51",
  1492 => x"848080d1",
  1493 => x"bb2d83ff",
  1494 => x"e0800879",
  1495 => x"0c848080",
  1496 => x"af890478",
  1497 => x"52941951",
  1498 => x"848080ab",
  1499 => x"982d83ff",
  1500 => x"e0800856",
  1501 => x"83ffe080",
  1502 => x"088f3878",
  1503 => x"51848080",
  1504 => x"aaf12d84",
  1505 => x"8080b0ef",
  1506 => x"0402a805",
  1507 => x"70558298",
  1508 => x"1a547908",
  1509 => x"5383ffe9",
  1510 => x"ec525684",
  1511 => x"8080d1ce",
  1512 => x"2d83ffe0",
  1513 => x"8008802e",
  1514 => x"81bb3875",
  1515 => x"51848080",
  1516 => x"a9882d83",
  1517 => x"ffe08008",
  1518 => x"802e81a9",
  1519 => x"388b5375",
  1520 => x"52849c19",
  1521 => x"51848080",
  1522 => x"ddd92d61",
  1523 => x"70882b87",
  1524 => x"fc808006",
  1525 => x"7072982b",
  1526 => x"0772882a",
  1527 => x"83fe8006",
  1528 => x"71077398",
  1529 => x"2a078c1d",
  1530 => x"0c515757",
  1531 => x"800b881a",
  1532 => x"0c02bc05",
  1533 => x"84808080",
  1534 => x"e02d7088",
  1535 => x"2b83fe80",
  1536 => x"0671882a",
  1537 => x"07028805",
  1538 => x"80c20584",
  1539 => x"808080e0",
  1540 => x"2d70882b",
  1541 => x"83fe8006",
  1542 => x"71882a07",
  1543 => x"72848080",
  1544 => x"2905841d",
  1545 => x"0c585158",
  1546 => x"ff0b88b0",
  1547 => x"1a0c800b",
  1548 => x"88b41a0c",
  1549 => x"800b901a",
  1550 => x"0cff0b84",
  1551 => x"a81a0cff",
  1552 => x"0b84ac1a",
  1553 => x"0c785283",
  1554 => x"ffe9ec51",
  1555 => x"848080c3",
  1556 => x"fb2d83ff",
  1557 => x"e9ec5184",
  1558 => x"80809481",
  1559 => x"2d785684",
  1560 => x"8080b0ef",
  1561 => x"04785184",
  1562 => x"8080aaf1",
  1563 => x"2d805675",
  1564 => x"83ffe080",
  1565 => x"0c0280c8",
  1566 => x"050d0402",
  1567 => x"d0050d7d",
  1568 => x"7f6283ff",
  1569 => x"e9ec0b84",
  1570 => x"808080f5",
  1571 => x"2d705672",
  1572 => x"555a5c56",
  1573 => x"59848080",
  1574 => x"e3842d83",
  1575 => x"ffe08008",
  1576 => x"83ffe080",
  1577 => x"08782976",
  1578 => x"71317c11",
  1579 => x"585d5758",
  1580 => x"76752785",
  1581 => x"38767b31",
  1582 => x"5a84a819",
  1583 => x"08567776",
  1584 => x"2e098106",
  1585 => x"8c3884ac",
  1586 => x"19085684",
  1587 => x"8080b2d9",
  1588 => x"0477802e",
  1589 => x"99388116",
  1590 => x"5577752e",
  1591 => x"0981068e",
  1592 => x"387584ac",
  1593 => x"1a085755",
  1594 => x"848080b1",
  1595 => x"f504800b",
  1596 => x"841a0857",
  1597 => x"55747827",
  1598 => x"80d03802",
  1599 => x"b005fc05",
  1600 => x"54745378",
  1601 => x"5283ffe9",
  1602 => x"ec518480",
  1603 => x"80c4832d",
  1604 => x"83ffe080",
  1605 => x"08a93875",
  1606 => x"5283ffe9",
  1607 => x"ec518480",
  1608 => x"8094ce2d",
  1609 => x"83ffe080",
  1610 => x"085c83ff",
  1611 => x"e0800854",
  1612 => x"74537852",
  1613 => x"83ffe9ec",
  1614 => x"51848080",
  1615 => x"c48b2d7b",
  1616 => x"81165656",
  1617 => x"848080b1",
  1618 => x"f50475ff",
  1619 => x"2e933875",
  1620 => x"84ac1a0c",
  1621 => x"7784a81a",
  1622 => x"0c75ff2e",
  1623 => x"09810689",
  1624 => x"38805584",
  1625 => x"8080b39b",
  1626 => x"04755283",
  1627 => x"ffe9ec51",
  1628 => x"848080cc",
  1629 => x"a62d7954",
  1630 => x"7f5383ff",
  1631 => x"e080081b",
  1632 => x"5283ffe9",
  1633 => x"ec518480",
  1634 => x"80ccfd2d",
  1635 => x"795583ff",
  1636 => x"e0800887",
  1637 => x"3883ffe0",
  1638 => x"80085574",
  1639 => x"83ffe080",
  1640 => x"0c02b005",
  1641 => x"0d0402f8",
  1642 => x"050d83ff",
  1643 => x"f2dc5184",
  1644 => x"8080a9b1",
  1645 => x"2d83fff2",
  1646 => x"d4518480",
  1647 => x"80a9b12d",
  1648 => x"83ffe9e4",
  1649 => x"5283fff2",
  1650 => x"dc518480",
  1651 => x"80a9fe2d",
  1652 => x"810b83ff",
  1653 => x"e1a00c02",
  1654 => x"88050d04",
  1655 => x"02fc050d",
  1656 => x"83ffeaa8",
  1657 => x"73717084",
  1658 => x"05530c74",
  1659 => x"710c5102",
  1660 => x"84050d04",
  1661 => x"02f4050d",
  1662 => x"83ffe1a0",
  1663 => x"08873884",
  1664 => x"8080b3a6",
  1665 => x"2d7483ff",
  1666 => x"eaa00c75",
  1667 => x"83ffeaa4",
  1668 => x"0c83ffe9",
  1669 => x"ec518480",
  1670 => x"80c4932d",
  1671 => x"83ffe080",
  1672 => x"085383ff",
  1673 => x"e0800880",
  1674 => x"2e993883",
  1675 => x"ffe08008",
  1676 => x"52848080",
  1677 => x"e7f85184",
  1678 => x"808082e3",
  1679 => x"2d848080",
  1680 => x"b4d00481",
  1681 => x"0b83ffe1",
  1682 => x"a40c83ff",
  1683 => x"e0800853",
  1684 => x"7283ffe0",
  1685 => x"800c028c",
  1686 => x"050d0402",
  1687 => x"f8050d83",
  1688 => x"ffe1a008",
  1689 => x"87388480",
  1690 => x"80b3a62d",
  1691 => x"83ffeaa8",
  1692 => x"08527180",
  1693 => x"2e833871",
  1694 => x"2d83ffe9",
  1695 => x"ec518480",
  1696 => x"8094812d",
  1697 => x"83ffeaac",
  1698 => x"08527180",
  1699 => x"2e833871",
  1700 => x"2d028805",
  1701 => x"0d0402e8",
  1702 => x"050d7779",
  1703 => x"56568054",
  1704 => x"83ffe1a0",
  1705 => x"08742e09",
  1706 => x"81068738",
  1707 => x"848080b3",
  1708 => x"a62d7352",
  1709 => x"83ffe1a4",
  1710 => x"08802e82",
  1711 => x"ff387581",
  1712 => x"05097077",
  1713 => x"07802576",
  1714 => x"81050970",
  1715 => x"78078025",
  1716 => x"72077752",
  1717 => x"52545153",
  1718 => x"7282e138",
  1719 => x"73538480",
  1720 => x"80b7b904",
  1721 => x"72157084",
  1722 => x"808080f5",
  1723 => x"2d515271",
  1724 => x"80d72e80",
  1725 => x"e8387180",
  1726 => x"d724ad38",
  1727 => x"7180c22e",
  1728 => x"81b03871",
  1729 => x"80c22494",
  1730 => x"3871ab2e",
  1731 => x"80e33871",
  1732 => x"80c12e80",
  1733 => x"d2388480",
  1734 => x"80b7b604",
  1735 => x"7180d22e",
  1736 => x"b2388480",
  1737 => x"80b7b604",
  1738 => x"7180e22e",
  1739 => x"81843871",
  1740 => x"80e2248d",
  1741 => x"387180e1",
  1742 => x"2ead3884",
  1743 => x"8080b7b6",
  1744 => x"047180f2",
  1745 => x"2e8d3871",
  1746 => x"80f72e91",
  1747 => x"38848080",
  1748 => x"b7b60473",
  1749 => x"81075484",
  1750 => x"8080b7b6",
  1751 => x"0473b207",
  1752 => x"54848080",
  1753 => x"b7b60473",
  1754 => x"a6075484",
  1755 => x"8080b7b6",
  1756 => x"04738106",
  1757 => x"5271802e",
  1758 => x"8b387382",
  1759 => x"07548480",
  1760 => x"80b7b604",
  1761 => x"73812a70",
  1762 => x"81065152",
  1763 => x"71802e8b",
  1764 => x"3873b107",
  1765 => x"54848080",
  1766 => x"b7b60473",
  1767 => x"822a7081",
  1768 => x"06515271",
  1769 => x"802e8f38",
  1770 => x"73a70754",
  1771 => x"848080b7",
  1772 => x"b6047388",
  1773 => x"07548113",
  1774 => x"53745184",
  1775 => x"8080d8ce",
  1776 => x"2d83ffe0",
  1777 => x"80087324",
  1778 => x"fe9a3880",
  1779 => x"7481d906",
  1780 => x"555383ff",
  1781 => x"eaa40873",
  1782 => x"2e098106",
  1783 => x"86387381",
  1784 => x"d9065483",
  1785 => x"ffeaa808",
  1786 => x"5271802e",
  1787 => x"8338712d",
  1788 => x"73810652",
  1789 => x"719a3873",
  1790 => x"852a7081",
  1791 => x"06515272",
  1792 => x"a2387180",
  1793 => x"2e983873",
  1794 => x"86065271",
  1795 => x"802e8f38",
  1796 => x"75518480",
  1797 => x"80ad832d",
  1798 => x"83ffe080",
  1799 => x"08537280",
  1800 => x"2e8b3873",
  1801 => x"88b81484",
  1802 => x"808081b7",
  1803 => x"2d83ffea",
  1804 => x"ac085271",
  1805 => x"802e8338",
  1806 => x"712d7252",
  1807 => x"7183ffe0",
  1808 => x"800c0298",
  1809 => x"050d0480",
  1810 => x"0b83ffe0",
  1811 => x"800c0402",
  1812 => x"f4050d74",
  1813 => x"5283ffe1",
  1814 => x"a0088738",
  1815 => x"848080b3",
  1816 => x"a62d7180",
  1817 => x"2e80da38",
  1818 => x"83ffeaa8",
  1819 => x"08537280",
  1820 => x"2e833872",
  1821 => x"2d901208",
  1822 => x"802e8638",
  1823 => x"800b9013",
  1824 => x"0c800b88",
  1825 => x"130c800b",
  1826 => x"8c130c80",
  1827 => x"0b84130c",
  1828 => x"ff0b88b0",
  1829 => x"130c800b",
  1830 => x"88b4130c",
  1831 => x"800b9013",
  1832 => x"0c715184",
  1833 => x"8080aaf1",
  1834 => x"2d83ffe9",
  1835 => x"ec518480",
  1836 => x"8094812d",
  1837 => x"83ffeaac",
  1838 => x"08527180",
  1839 => x"2e833871",
  1840 => x"2d028c05",
  1841 => x"0d0402d0",
  1842 => x"050d7d61",
  1843 => x"6062295a",
  1844 => x"5a5c805b",
  1845 => x"83ffe1a0",
  1846 => x"087b2e09",
  1847 => x"81068738",
  1848 => x"848080b3",
  1849 => x"a62d7b81",
  1850 => x"0509707d",
  1851 => x"0780257a",
  1852 => x"81050970",
  1853 => x"7c078025",
  1854 => x"72075257",
  1855 => x"5156ff5a",
  1856 => x"7581f238",
  1857 => x"88b81984",
  1858 => x"808080f5",
  1859 => x"2d810655",
  1860 => x"74802e81",
  1861 => x"e0387a5a",
  1862 => x"77802e81",
  1863 => x"d8388819",
  1864 => x"088c1a08",
  1865 => x"5856ff5a",
  1866 => x"75772781",
  1867 => x"c8387716",
  1868 => x"55767527",
  1869 => x"85387676",
  1870 => x"31587589",
  1871 => x"2a7683ff",
  1872 => x"065b5580",
  1873 => x"782581ab",
  1874 => x"387980c4",
  1875 => x"38777b31",
  1876 => x"5683ff76",
  1877 => x"25ba3875",
  1878 => x"80258538",
  1879 => x"83ff1656",
  1880 => x"75892c54",
  1881 => x"7a1c5374",
  1882 => x"52785184",
  1883 => x"8080b0fb",
  1884 => x"2d83ffe0",
  1885 => x"8008802e",
  1886 => x"80f93883",
  1887 => x"ffe08008",
  1888 => x"892b83ff",
  1889 => x"e0800816",
  1890 => x"56578480",
  1891 => x"80bbe304",
  1892 => x"88b01908",
  1893 => x"752ea638",
  1894 => x"815484b0",
  1895 => x"19537452",
  1896 => x"78518480",
  1897 => x"80b0fb2d",
  1898 => x"83ffe080",
  1899 => x"08802e80",
  1900 => x"c2387488",
  1901 => x"b01a0c80",
  1902 => x"0b88b41a",
  1903 => x"0c84807a",
  1904 => x"31787c31",
  1905 => x"57577577",
  1906 => x"25833875",
  1907 => x"57765379",
  1908 => x"1984b005",
  1909 => x"527a1c51",
  1910 => x"848080dd",
  1911 => x"d92d8115",
  1912 => x"55805a76",
  1913 => x"1b881a08",
  1914 => x"18881b0c",
  1915 => x"5b777b24",
  1916 => x"fed7387a",
  1917 => x"5a7983ff",
  1918 => x"e0800c02",
  1919 => x"b0050d04",
  1920 => x"02e8050d",
  1921 => x"80029805",
  1922 => x"84808081",
  1923 => x"b72d7754",
  1924 => x"81538152",
  1925 => x"029805fc",
  1926 => x"05518480",
  1927 => x"80b9c62d",
  1928 => x"83ffe080",
  1929 => x"085583ff",
  1930 => x"e0800881",
  1931 => x"2e098106",
  1932 => x"8b380294",
  1933 => x"05848080",
  1934 => x"80f52d55",
  1935 => x"7483ffe0",
  1936 => x"800c0298",
  1937 => x"050d0402",
  1938 => x"e8050d77",
  1939 => x"797b5853",
  1940 => x"55805372",
  1941 => x"722580d4",
  1942 => x"38ff1254",
  1943 => x"72742580",
  1944 => x"cb387551",
  1945 => x"848080bc",
  1946 => x"802d800b",
  1947 => x"83ffe080",
  1948 => x"0824a138",
  1949 => x"74135283",
  1950 => x"ffe08008",
  1951 => x"72848080",
  1952 => x"81b72d81",
  1953 => x"135383ff",
  1954 => x"e080088a",
  1955 => x"2e863873",
  1956 => x"7324cf38",
  1957 => x"80732594",
  1958 => x"38721552",
  1959 => x"80728480",
  1960 => x"8081b72d",
  1961 => x"74528480",
  1962 => x"80bdae04",
  1963 => x"80527183",
  1964 => x"ffe0800c",
  1965 => x"0298050d",
  1966 => x"0402e805",
  1967 => x"0d77797b",
  1968 => x"585454ff",
  1969 => x"5583ffe1",
  1970 => x"a0088738",
  1971 => x"848080b3",
  1972 => x"a62d7452",
  1973 => x"73802e81",
  1974 => x"bc387582",
  1975 => x"32708105",
  1976 => x"09707207",
  1977 => x"80255152",
  1978 => x"5272802e",
  1979 => x"87387452",
  1980 => x"7081a238",
  1981 => x"83ffeaa8",
  1982 => x"08517080",
  1983 => x"2e833870",
  1984 => x"2dff0b88",
  1985 => x"b0150c80",
  1986 => x"0b88b415",
  1987 => x"0c759a38",
  1988 => x"7288150c",
  1989 => x"8c140851",
  1990 => x"70732785",
  1991 => x"38708815",
  1992 => x"0c755584",
  1993 => x"8080bf86",
  1994 => x"0475812e",
  1995 => x"09810680",
  1996 => x"c5388814",
  1997 => x"08518073",
  1998 => x"249b3872",
  1999 => x"11708816",
  2000 => x"0c8c1508",
  2001 => x"53517171",
  2002 => x"27ba3871",
  2003 => x"88150c84",
  2004 => x"8080bf84",
  2005 => x"04728105",
  2006 => x"09537073",
  2007 => x"278c3880",
  2008 => x"0b88150c",
  2009 => x"848080bf",
  2010 => x"84047073",
  2011 => x"3188150c",
  2012 => x"848080bf",
  2013 => x"84047582",
  2014 => x"2e098106",
  2015 => x"89388c14",
  2016 => x"0888150c",
  2017 => x"805583ff",
  2018 => x"eaac0851",
  2019 => x"70802e83",
  2020 => x"38702d74",
  2021 => x"527183ff",
  2022 => x"e0800c02",
  2023 => x"98050d04",
  2024 => x"02f8050d",
  2025 => x"7352ff51",
  2026 => x"71802ea4",
  2027 => x"3883ffea",
  2028 => x"a8085170",
  2029 => x"802e8338",
  2030 => x"702d7488",
  2031 => x"1308710c",
  2032 => x"5183ffea",
  2033 => x"ac085170",
  2034 => x"802e8338",
  2035 => x"702d8051",
  2036 => x"7083ffe0",
  2037 => x"800c0288",
  2038 => x"050d0402",
  2039 => x"f0050d80",
  2040 => x"54029005",
  2041 => x"fc055275",
  2042 => x"51848080",
  2043 => x"bfa02d73",
  2044 => x"83ffe080",
  2045 => x"0c029005",
  2046 => x"0d0402f8",
  2047 => x"050d7352",
  2048 => x"ff517180",
  2049 => x"2eb13883",
  2050 => x"ffeaa808",
  2051 => x"5170802e",
  2052 => x"8338702d",
  2053 => x"8812088c",
  2054 => x"13083270",
  2055 => x"81050970",
  2056 => x"72079f2a",
  2057 => x"ff1183ff",
  2058 => x"eaac0854",
  2059 => x"51515252",
  2060 => x"71802e83",
  2061 => x"38712d70",
  2062 => x"83ffe080",
  2063 => x"0c028805",
  2064 => x"0d04800b",
  2065 => x"83ffe080",
  2066 => x"0c0402e4",
  2067 => x"050d787a",
  2068 => x"5755ff57",
  2069 => x"83ffe1a0",
  2070 => x"08873884",
  2071 => x"8080b3a6",
  2072 => x"2d83ffea",
  2073 => x"a8085473",
  2074 => x"802e8338",
  2075 => x"732d7451",
  2076 => x"84808099",
  2077 => x"cb2d83ff",
  2078 => x"e08008ff",
  2079 => x"2e098106",
  2080 => x"983883ff",
  2081 => x"e9ec5184",
  2082 => x"8080d1bb",
  2083 => x"2d83ffe0",
  2084 => x"80085784",
  2085 => x"8080c1b0",
  2086 => x"04029c05",
  2087 => x"fc055274",
  2088 => x"51848080",
  2089 => x"ab982d83",
  2090 => x"ffe08008",
  2091 => x"802e9038",
  2092 => x"76537552",
  2093 => x"83ffe9ec",
  2094 => x"51848080",
  2095 => x"d49d2d83",
  2096 => x"ffeaac08",
  2097 => x"5473802e",
  2098 => x"8338732d",
  2099 => x"755476ff",
  2100 => x"2e098106",
  2101 => x"83388054",
  2102 => x"7383ffe0",
  2103 => x"800c029c",
  2104 => x"050d0402",
  2105 => x"ec050d83",
  2106 => x"ffe1a008",
  2107 => x"87388480",
  2108 => x"80b3a62d",
  2109 => x"83ffeaa8",
  2110 => x"08547380",
  2111 => x"2e833873",
  2112 => x"2d775376",
  2113 => x"5283ffe9",
  2114 => x"ec518480",
  2115 => x"80d4b92d",
  2116 => x"83ffe080",
  2117 => x"0883ffea",
  2118 => x"ac085555",
  2119 => x"73802e83",
  2120 => x"38732d74",
  2121 => x"83ffe080",
  2122 => x"0c029405",
  2123 => x"0d0402fd",
  2124 => x"cc050d83",
  2125 => x"ffe1a008",
  2126 => x"87388480",
  2127 => x"80b3a62d",
  2128 => x"83ffeaa8",
  2129 => x"08547380",
  2130 => x"2e833873",
  2131 => x"2d0282a8",
  2132 => x"05705302",
  2133 => x"82bc0508",
  2134 => x"52568480",
  2135 => x"80c0ca2d",
  2136 => x"83ffe080",
  2137 => x"08802e80",
  2138 => x"d5388480",
  2139 => x"80c3a804",
  2140 => x"02829c05",
  2141 => x"84808080",
  2142 => x"f52d5473",
  2143 => x"802e9538",
  2144 => x"74528480",
  2145 => x"80e8ac51",
  2146 => x"84808082",
  2147 => x"e32d8480",
  2148 => x"80c3a804",
  2149 => x"0282a405",
  2150 => x"08537452",
  2151 => x"848080e8",
  2152 => x"b8518480",
  2153 => x"8082e32d",
  2154 => x"02980570",
  2155 => x"53765255",
  2156 => x"848080c1",
  2157 => x"e32d83ff",
  2158 => x"e08008ff",
  2159 => x"b33883ff",
  2160 => x"eaac0854",
  2161 => x"73802e83",
  2162 => x"38732d02",
  2163 => x"82b4050d",
  2164 => x"0402e405",
  2165 => x"0d8002a0",
  2166 => x"05f40553",
  2167 => x"79525384",
  2168 => x"8080c0ca",
  2169 => x"2d83ffe0",
  2170 => x"8008732e",
  2171 => x"83388153",
  2172 => x"7283ffe0",
  2173 => x"800c029c",
  2174 => x"050d0481",
  2175 => x"0b83ffe0",
  2176 => x"800c0480",
  2177 => x"0b83ffe0",
  2178 => x"800c0481",
  2179 => x"0b83ffe0",
  2180 => x"800c0402",
  2181 => x"ffb8050d",
  2182 => x"63578058",
  2183 => x"ff0b84c4",
  2184 => x"180c7784",
  2185 => x"c8180c77",
  2186 => x"a4180c76",
  2187 => x"51848080",
  2188 => x"90f92db4",
  2189 => x"170854ff",
  2190 => x"5573782e",
  2191 => x"87dc3881",
  2192 => x"5380c417",
  2193 => x"70537852",
  2194 => x"59732d83",
  2195 => x"ffe08008",
  2196 => x"782e87c6",
  2197 => x"3884c217",
  2198 => x"84808080",
  2199 => x"e02d54fd",
  2200 => x"557381ab",
  2201 => x"aa2e0981",
  2202 => x"0687af38",
  2203 => x"84c31784",
  2204 => x"808080f5",
  2205 => x"2d84c218",
  2206 => x"84808080",
  2207 => x"f52d7182",
  2208 => x"80290555",
  2209 => x"55fc5573",
  2210 => x"82d4d52e",
  2211 => x"09810687",
  2212 => x"89388486",
  2213 => x"17848080",
  2214 => x"80f52d70",
  2215 => x"81ff0655",
  2216 => x"56738f26",
  2217 => x"a0388174",
  2218 => x"2b7083b0",
  2219 => x"e0065555",
  2220 => x"73782e09",
  2221 => x"81069938",
  2222 => x"74810654",
  2223 => x"73782e09",
  2224 => x"810680d0",
  2225 => x"387581ff",
  2226 => x"06547386",
  2227 => x"2680c538",
  2228 => x"848d1784",
  2229 => x"808080f5",
  2230 => x"2d848c18",
  2231 => x"84808080",
  2232 => x"f52d7181",
  2233 => x"800a2971",
  2234 => x"84808029",
  2235 => x"05848b1a",
  2236 => x"84808080",
  2237 => x"f52d7082",
  2238 => x"80291284",
  2239 => x"8a1c8480",
  2240 => x"8080f52d",
  2241 => x"5574059c",
  2242 => x"1c0c5956",
  2243 => x"56588480",
  2244 => x"80c69804",
  2245 => x"779c180c",
  2246 => x"81537852",
  2247 => x"9c170851",
  2248 => x"b4170854",
  2249 => x"732dff55",
  2250 => x"83ffe080",
  2251 => x"08802e85",
  2252 => x"e93880d0",
  2253 => x"17848080",
  2254 => x"80f52d80",
  2255 => x"cf188480",
  2256 => x"8080f52d",
  2257 => x"7072882b",
  2258 => x"0756415f",
  2259 => x"fe557384",
  2260 => x"802e0981",
  2261 => x"0685c338",
  2262 => x"80d11784",
  2263 => x"808080f5",
  2264 => x"2d778480",
  2265 => x"8081b72d",
  2266 => x"80d31784",
  2267 => x"808080f5",
  2268 => x"2d80d218",
  2269 => x"84808080",
  2270 => x"f52d7072",
  2271 => x"882b0780",
  2272 => x"d41a8480",
  2273 => x"8080f52d",
  2274 => x"7081ff06",
  2275 => x"80d61c84",
  2276 => x"808080f5",
  2277 => x"2d80d51d",
  2278 => x"84808080",
  2279 => x"f52d7072",
  2280 => x"882b075b",
  2281 => x"415f5a41",
  2282 => x"5b434173",
  2283 => x"a8188480",
  2284 => x"80818a2d",
  2285 => x"80db1784",
  2286 => x"808080f5",
  2287 => x"2d80da18",
  2288 => x"84808080",
  2289 => x"f52d7072",
  2290 => x"882b0756",
  2291 => x"5e5c7380",
  2292 => x"2e8b3873",
  2293 => x"a0180c84",
  2294 => x"8080c89b",
  2295 => x"0480eb17",
  2296 => x"84808080",
  2297 => x"f52d80ea",
  2298 => x"18848080",
  2299 => x"80f52d71",
  2300 => x"81800a29",
  2301 => x"71848080",
  2302 => x"290580e9",
  2303 => x"1a848080",
  2304 => x"80f52d70",
  2305 => x"82802912",
  2306 => x"80e81c84",
  2307 => x"808080f5",
  2308 => x"2d547305",
  2309 => x"a01c0c53",
  2310 => x"56595580",
  2311 => x"f3178480",
  2312 => x"8080f52d",
  2313 => x"80f21884",
  2314 => x"808080f5",
  2315 => x"2d718180",
  2316 => x"0a297184",
  2317 => x"80802905",
  2318 => x"80f11a84",
  2319 => x"808080f5",
  2320 => x"2d708280",
  2321 => x"291280f0",
  2322 => x"1c848080",
  2323 => x"80f52d54",
  2324 => x"7305881c",
  2325 => x"0c80f51b",
  2326 => x"84808080",
  2327 => x"f52d80f4",
  2328 => x"1c848080",
  2329 => x"80f52d71",
  2330 => x"82802905",
  2331 => x"53515356",
  2332 => x"59557398",
  2333 => x"18848080",
  2334 => x"818a2d75",
  2335 => x"a0180829",
  2336 => x"701a8c19",
  2337 => x"0ca81884",
  2338 => x"808080e0",
  2339 => x"2d70852b",
  2340 => x"83ff1152",
  2341 => x"58555873",
  2342 => x"80258538",
  2343 => x"87fe1654",
  2344 => x"73892a90",
  2345 => x"180c9c17",
  2346 => x"08197094",
  2347 => x"190c7805",
  2348 => x"84180c84",
  2349 => x"c3178480",
  2350 => x"8080f52d",
  2351 => x"84c21884",
  2352 => x"808080f5",
  2353 => x"2d718280",
  2354 => x"29055555",
  2355 => x"fd557382",
  2356 => x"d4d52e09",
  2357 => x"810682c2",
  2358 => x"3879882b",
  2359 => x"83fe8006",
  2360 => x"7b81ff06",
  2361 => x"7012852b",
  2362 => x"61882b83",
  2363 => x"fe800663",
  2364 => x"81ff0671",
  2365 => x"05705751",
  2366 => x"527105ff",
  2367 => x"05535556",
  2368 => x"848080e2",
  2369 => x"b12d83ff",
  2370 => x"e080087c",
  2371 => x"882b83fe",
  2372 => x"80067e81",
  2373 => x"ff067105",
  2374 => x"705c5155",
  2375 => x"5a73bd38",
  2376 => x"80eb1784",
  2377 => x"808080f5",
  2378 => x"2d80ea18",
  2379 => x"84808080",
  2380 => x"f52d7181",
  2381 => x"800a2971",
  2382 => x"84808029",
  2383 => x"0580e91a",
  2384 => x"84808080",
  2385 => x"f52d7082",
  2386 => x"80291280",
  2387 => x"e81c8480",
  2388 => x"8080f52d",
  2389 => x"5574055d",
  2390 => x"59565658",
  2391 => x"80d81784",
  2392 => x"808080f5",
  2393 => x"2d80d718",
  2394 => x"84808080",
  2395 => x"f52d7182",
  2396 => x"80290570",
  2397 => x"5a555573",
  2398 => x"bd3880e7",
  2399 => x"17848080",
  2400 => x"80f52d80",
  2401 => x"e6188480",
  2402 => x"8080f52d",
  2403 => x"7181800a",
  2404 => x"29718480",
  2405 => x"80290580",
  2406 => x"e51a8480",
  2407 => x"8080f52d",
  2408 => x"70828029",
  2409 => x"1280e41c",
  2410 => x"84808080",
  2411 => x"f52d5473",
  2412 => x"05545956",
  2413 => x"56586088",
  2414 => x"2b83fe80",
  2415 => x"066281ff",
  2416 => x"067f81ff",
  2417 => x"06577105",
  2418 => x"767b2905",
  2419 => x"7971317c",
  2420 => x"31798480",
  2421 => x"8080f52d",
  2422 => x"52585154",
  2423 => x"fb557380",
  2424 => x"2eb83873",
  2425 => x"52755184",
  2426 => x"8080e384",
  2427 => x"2d9ff40b",
  2428 => x"83ffe080",
  2429 => x"0827a338",
  2430 => x"83ffe080",
  2431 => x"0883fff4",
  2432 => x"26913880",
  2433 => x"0b88180c",
  2434 => x"800bb018",
  2435 => x"0c848080",
  2436 => x"cc980481",
  2437 => x"0bb0180c",
  2438 => x"80557483",
  2439 => x"ffe0800c",
  2440 => x"0280c805",
  2441 => x"0d0402e8",
  2442 => x"050d7779",
  2443 => x"5755b015",
  2444 => x"08af38a8",
  2445 => x"15848080",
  2446 => x"80e02d53",
  2447 => x"72802584",
  2448 => x"388f1353",
  2449 => x"72842a84",
  2450 => x"16080575",
  2451 => x"84808080",
  2452 => x"f52dfe18",
  2453 => x"71297205",
  2454 => x"52565484",
  2455 => x"8080ccf2",
  2456 => x"04748480",
  2457 => x"8080f52d",
  2458 => x"fe177129",
  2459 => x"84170805",
  2460 => x"51547383",
  2461 => x"ffe0800c",
  2462 => x"0298050d",
  2463 => x"0402f005",
  2464 => x"0d785377",
  2465 => x"52765175",
  2466 => x"b4110851",
  2467 => x"54732d02",
  2468 => x"90050d04",
  2469 => x"02f0050d",
  2470 => x"78537752",
  2471 => x"765175b8",
  2472 => x"11085154",
  2473 => x"732d0290",
  2474 => x"050d0402",
  2475 => x"d4050d7c",
  2476 => x"7e60625e",
  2477 => x"5c565780",
  2478 => x"705559b0",
  2479 => x"1708792e",
  2480 => x"09810683",
  2481 => x"38815478",
  2482 => x"5874a138",
  2483 => x"73587380",
  2484 => x"2e9a3878",
  2485 => x"55799018",
  2486 => x"082781a0",
  2487 => x"389c1708",
  2488 => x"8c180805",
  2489 => x"1a548480",
  2490 => x"80ceca04",
  2491 => x"74778480",
  2492 => x"8080f52d",
  2493 => x"70547b53",
  2494 => x"55568480",
  2495 => x"80e3842d",
  2496 => x"83ffe080",
  2497 => x"0874297a",
  2498 => x"71315a54",
  2499 => x"7783ffe0",
  2500 => x"8008279d",
  2501 => x"3883ffe0",
  2502 => x"80085475",
  2503 => x"52765184",
  2504 => x"808094ce",
  2505 => x"2d83ffe0",
  2506 => x"8008ff15",
  2507 => x"555673eb",
  2508 => x"38805575",
  2509 => x"ff2e80c4",
  2510 => x"38755276",
  2511 => x"51848080",
  2512 => x"cca62d83",
  2513 => x"ffe08008",
  2514 => x"19547a80",
  2515 => x"2e8b3881",
  2516 => x"537a5284",
  2517 => x"8080ceee",
  2518 => x"04815573",
  2519 => x"84c41808",
  2520 => x"2e9a3873",
  2521 => x"84c4180c",
  2522 => x"745380c4",
  2523 => x"17527351",
  2524 => x"b4170854",
  2525 => x"732d83ff",
  2526 => x"e0800855",
  2527 => x"7483ffe0",
  2528 => x"800c02ac",
  2529 => x"050d0402",
  2530 => x"d8050d7b",
  2531 => x"7d7f61b0",
  2532 => x"14087081",
  2533 => x"0509b016",
  2534 => x"08710770",
  2535 => x"09709f2a",
  2536 => x"51515151",
  2537 => x"585c5c59",
  2538 => x"5677bf38",
  2539 => x"81707506",
  2540 => x"55577380",
  2541 => x"2eb43877",
  2542 => x"54799017",
  2543 => x"082780f4",
  2544 => x"389c1608",
  2545 => x"8c170805",
  2546 => x"1ab41708",
  2547 => x"56547880",
  2548 => x"2e8b3876",
  2549 => x"53785284",
  2550 => x"8080d0aa",
  2551 => x"047384c4",
  2552 => x"170c7653",
  2553 => x"848080d0",
  2554 => x"a604b416",
  2555 => x"08557880",
  2556 => x"2e9c3877",
  2557 => x"52755184",
  2558 => x"8080cca6",
  2559 => x"2d815378",
  2560 => x"5283ffe0",
  2561 => x"80081a51",
  2562 => x"848080d0",
  2563 => x"ac047752",
  2564 => x"75518480",
  2565 => x"80cca62d",
  2566 => x"83ffe080",
  2567 => x"081a7084",
  2568 => x"c4180c54",
  2569 => x"815380c4",
  2570 => x"16527351",
  2571 => x"742d83ff",
  2572 => x"e0800854",
  2573 => x"7383ffe0",
  2574 => x"800c02a8",
  2575 => x"050d0402",
  2576 => x"f0050d75",
  2577 => x"848080e8",
  2578 => x"c8525484",
  2579 => x"808082e3",
  2580 => x"2d848080",
  2581 => x"e8d853b0",
  2582 => x"1408812e",
  2583 => x"87388480",
  2584 => x"80e8e053",
  2585 => x"72528480",
  2586 => x"80e8e851",
  2587 => x"84808082",
  2588 => x"e32d8814",
  2589 => x"08528480",
  2590 => x"80e8f451",
  2591 => x"84808082",
  2592 => x"e32d9414",
  2593 => x"08528480",
  2594 => x"80e99451",
  2595 => x"84808082",
  2596 => x"e32d8414",
  2597 => x"08528480",
  2598 => x"80e9ac51",
  2599 => x"84808082",
  2600 => x"e32d7384",
  2601 => x"808080f5",
  2602 => x"2d528480",
  2603 => x"80e9c851",
  2604 => x"84808082",
  2605 => x"e32d0290",
  2606 => x"050d0402",
  2607 => x"fc050d72",
  2608 => x"88110883",
  2609 => x"ffe0800c",
  2610 => x"51028405",
  2611 => x"0d0402ff",
  2612 => x"ac050d66",
  2613 => x"686a4141",
  2614 => x"5e805d81",
  2615 => x"520280d4",
  2616 => x"05ec0551",
  2617 => x"848080a7",
  2618 => x"df2d8054",
  2619 => x"7c53811d",
  2620 => x"60537e52",
  2621 => x"5d848080",
  2622 => x"cdab2d83",
  2623 => x"ffe08008",
  2624 => x"802e828b",
  2625 => x"38805b7a",
  2626 => x"a0291e80",
  2627 => x"c4057052",
  2628 => x"58848080",
  2629 => x"a89b2d83",
  2630 => x"ffe08008",
  2631 => x"802e81db",
  2632 => x"380280c4",
  2633 => x"05598d53",
  2634 => x"80527851",
  2635 => x"848080e0",
  2636 => x"cc2d8057",
  2637 => x"76197719",
  2638 => x"57557584",
  2639 => x"808080f5",
  2640 => x"2d758480",
  2641 => x"8081b72d",
  2642 => x"81177081",
  2643 => x"ff065855",
  2644 => x"877727e0",
  2645 => x"38805a88",
  2646 => x"02840580",
  2647 => x"c5055d57",
  2648 => x"761c7719",
  2649 => x"56567484",
  2650 => x"808080f5",
  2651 => x"2d768480",
  2652 => x"8081b72d",
  2653 => x"74848080",
  2654 => x"80f52d55",
  2655 => x"74a02e83",
  2656 => x"38815a81",
  2657 => x"177081ff",
  2658 => x"0658558a",
  2659 => x"7727d138",
  2660 => x"79802ea2",
  2661 => x"380280c4",
  2662 => x"05848080",
  2663 => x"80f52d55",
  2664 => x"74ae2e92",
  2665 => x"38ae0280",
  2666 => x"d0058480",
  2667 => x"8081b72d",
  2668 => x"848080d3",
  2669 => x"c104a002",
  2670 => x"80d00584",
  2671 => x"808081b7",
  2672 => x"2d7e5278",
  2673 => x"51848080",
  2674 => x"a09e2d83",
  2675 => x"ffe08008",
  2676 => x"802e9538",
  2677 => x"a0537752",
  2678 => x"69518480",
  2679 => x"80ddd92d",
  2680 => x"81558480",
  2681 => x"80d49104",
  2682 => x"83ffe080",
  2683 => x"08520280",
  2684 => x"d405ec05",
  2685 => x"51848080",
  2686 => x"a7df2d81",
  2687 => x"1b7081ff",
  2688 => x"065c558f",
  2689 => x"7b27fdff",
  2690 => x"38848080",
  2691 => x"d1ea0480",
  2692 => x"557483ff",
  2693 => x"e0800c02",
  2694 => x"80d4050d",
  2695 => x"0402fc05",
  2696 => x"0d737584",
  2697 => x"120c5180",
  2698 => x"710c800b",
  2699 => x"88128480",
  2700 => x"8081b72d",
  2701 => x"0284050d",
  2702 => x"0402ffb4",
  2703 => x"050d6466",
  2704 => x"68405b56",
  2705 => x"80520280",
  2706 => x"cc05ec05",
  2707 => x"51848080",
  2708 => x"a7df2d80",
  2709 => x"54790853",
  2710 => x"841a0852",
  2711 => x"75518480",
  2712 => x"80cdab2d",
  2713 => x"83ffe080",
  2714 => x"08802e83",
  2715 => x"d338881a",
  2716 => x"84808080",
  2717 => x"f52d5978",
  2718 => x"8f2683ae",
  2719 => x"3878a029",
  2720 => x"1680c405",
  2721 => x"70525884",
  2722 => x"8080a89b",
  2723 => x"2d83ffe0",
  2724 => x"8008802e",
  2725 => x"83863880",
  2726 => x"520280cc",
  2727 => x"05ec0551",
  2728 => x"848080a7",
  2729 => x"df2d02bc",
  2730 => x"055b8d53",
  2731 => x"80527a51",
  2732 => x"848080e0",
  2733 => x"cc2d8057",
  2734 => x"761b7719",
  2735 => x"57557584",
  2736 => x"808080f5",
  2737 => x"2d758480",
  2738 => x"8081b72d",
  2739 => x"81177081",
  2740 => x"ff065855",
  2741 => x"877727e0",
  2742 => x"38805c88",
  2743 => x"028405bd",
  2744 => x"055e5776",
  2745 => x"1d771956",
  2746 => x"56748480",
  2747 => x"8080f52d",
  2748 => x"76848080",
  2749 => x"81b72d74",
  2750 => x"84808080",
  2751 => x"f52d5574",
  2752 => x"a02e8338",
  2753 => x"815c8117",
  2754 => x"7081ff06",
  2755 => x"58558a77",
  2756 => x"27d1387b",
  2757 => x"802ea138",
  2758 => x"02bc0584",
  2759 => x"808080f5",
  2760 => x"2d5574ae",
  2761 => x"2e9238ae",
  2762 => x"0280c805",
  2763 => x"84808081",
  2764 => x"b72d8480",
  2765 => x"80d6c304",
  2766 => x"a00280c8",
  2767 => x"05848080",
  2768 => x"81b72d7a",
  2769 => x"527d5184",
  2770 => x"8080a3d6",
  2771 => x"2d775184",
  2772 => x"8080a8df",
  2773 => x"2d83ffe0",
  2774 => x"8008802e",
  2775 => x"9238810b",
  2776 => x"82841f84",
  2777 => x"808081b7",
  2778 => x"2d848080",
  2779 => x"d6fd0483",
  2780 => x"ffe08008",
  2781 => x"82841f84",
  2782 => x"808081b7",
  2783 => x"2d9c1884",
  2784 => x"808080f5",
  2785 => x"2d9d1984",
  2786 => x"808080f5",
  2787 => x"2d71982b",
  2788 => x"71902b07",
  2789 => x"9e1b8480",
  2790 => x"8080f52d",
  2791 => x"70882b72",
  2792 => x"079f1d84",
  2793 => x"808080f5",
  2794 => x"2d710770",
  2795 => x"882b87fc",
  2796 => x"80800670",
  2797 => x"72982b07",
  2798 => x"72882a83",
  2799 => x"fe800671",
  2800 => x"0773982a",
  2801 => x"0766828c",
  2802 => x"050c5153",
  2803 => x"51525957",
  2804 => x"951a8480",
  2805 => x"8080f52d",
  2806 => x"941b8480",
  2807 => x"8080f52d",
  2808 => x"71982b71",
  2809 => x"902b079b",
  2810 => x"1d848080",
  2811 => x"80f52d9a",
  2812 => x"1e848080",
  2813 => x"80f52d71",
  2814 => x"882b0772",
  2815 => x"07648288",
  2816 => x"050c811f",
  2817 => x"53555a58",
  2818 => x"515c5774",
  2819 => x"881b8480",
  2820 => x"8081b72d",
  2821 => x"81558480",
  2822 => x"80d8c204",
  2823 => x"81197081",
  2824 => x"ff065a55",
  2825 => x"848080d4",
  2826 => x"f7047908",
  2827 => x"81057a0c",
  2828 => x"800b881b",
  2829 => x"84808081",
  2830 => x"b72d8480",
  2831 => x"80d4d304",
  2832 => x"80557483",
  2833 => x"ffe0800c",
  2834 => x"0280cc05",
  2835 => x"0d0402f4",
  2836 => x"050d7452",
  2837 => x"80727081",
  2838 => x"05548480",
  2839 => x"8080f52d",
  2840 => x"52537073",
  2841 => x"2e933881",
  2842 => x"13727081",
  2843 => x"05548480",
  2844 => x"8080f52d",
  2845 => x"525370ef",
  2846 => x"387283ff",
  2847 => x"e0800c02",
  2848 => x"8c050d04",
  2849 => x"02f0050d",
  2850 => x"75777156",
  2851 => x"54527270",
  2852 => x"81055484",
  2853 => x"808080f5",
  2854 => x"2d517072",
  2855 => x"70810554",
  2856 => x"84808081",
  2857 => x"b72d70e6",
  2858 => x"387383ff",
  2859 => x"e0800c02",
  2860 => x"90050d04",
  2861 => x"02e4050d",
  2862 => x"787a7c72",
  2863 => x"5a545553",
  2864 => x"848080d9",
  2865 => x"d5048114",
  2866 => x"54747370",
  2867 => x"81055584",
  2868 => x"808081b7",
  2869 => x"2d807484",
  2870 => x"808080f5",
  2871 => x"2d7081ff",
  2872 => x"06535656",
  2873 => x"70762e83",
  2874 => x"38815671",
  2875 => x"81050970",
  2876 => x"73079f2a",
  2877 => x"707806ff",
  2878 => x"15555151",
  2879 => x"5170c738",
  2880 => x"71ff2e96",
  2881 => x"38807370",
  2882 => x"81055584",
  2883 => x"808081b7",
  2884 => x"2dff1252",
  2885 => x"848080da",
  2886 => x"80047683",
  2887 => x"ffe0800c",
  2888 => x"029c050d",
  2889 => x"0402f005",
  2890 => x"0d757771",
  2891 => x"56545271",
  2892 => x"70810553",
  2893 => x"84808080",
  2894 => x"f52d5170",
  2895 => x"f2387270",
  2896 => x"81055484",
  2897 => x"808080f5",
  2898 => x"2d517072",
  2899 => x"70810554",
  2900 => x"84808081",
  2901 => x"b72d70e6",
  2902 => x"387383ff",
  2903 => x"e0800c02",
  2904 => x"90050d04",
  2905 => x"02ec050d",
  2906 => x"76787a72",
  2907 => x"58555552",
  2908 => x"71708105",
  2909 => x"53848080",
  2910 => x"80f52d51",
  2911 => x"70f23884",
  2912 => x"8080db93",
  2913 => x"04ff1353",
  2914 => x"72ff2e9a",
  2915 => x"38811281",
  2916 => x"15555273",
  2917 => x"84808080",
  2918 => x"f52d5170",
  2919 => x"72848080",
  2920 => x"81b72d70",
  2921 => x"e0388072",
  2922 => x"84808081",
  2923 => x"b72d7483",
  2924 => x"ffe0800c",
  2925 => x"0294050d",
  2926 => x"0402f005",
  2927 => x"0d757752",
  2928 => x"52848080",
  2929 => x"dbdd0470",
  2930 => x"84808080",
  2931 => x"f52d5472",
  2932 => x"742e0981",
  2933 => x"06923881",
  2934 => x"12811252",
  2935 => x"52718480",
  2936 => x"8080f52d",
  2937 => x"5372e038",
  2938 => x"71848080",
  2939 => x"80f52d71",
  2940 => x"84808080",
  2941 => x"f52d7171",
  2942 => x"3183ffe0",
  2943 => x"800c5252",
  2944 => x"0290050d",
  2945 => x"0402ec05",
  2946 => x"0d76787a",
  2947 => x"70555354",
  2948 => x"5470802e",
  2949 => x"80c33884",
  2950 => x"8080dcab",
  2951 => x"04ff1151",
  2952 => x"70802ea1",
  2953 => x"38811481",
  2954 => x"14545473",
  2955 => x"84808080",
  2956 => x"f52d5271",
  2957 => x"802e8e38",
  2958 => x"72848080",
  2959 => x"80f52d55",
  2960 => x"71752ed9",
  2961 => x"38738480",
  2962 => x"8080f52d",
  2963 => x"73848080",
  2964 => x"80f52d71",
  2965 => x"71315454",
  2966 => x"547183ff",
  2967 => x"e0800c02",
  2968 => x"94050d04",
  2969 => x"02f4050d",
  2970 => x"74765451",
  2971 => x"848080dc",
  2972 => x"fa047173",
  2973 => x"2e8f3881",
  2974 => x"11517084",
  2975 => x"808080f5",
  2976 => x"2d5271ee",
  2977 => x"387083ff",
  2978 => x"e0800c02",
  2979 => x"8c050d04",
  2980 => x"02ec050d",
  2981 => x"76785653",
  2982 => x"80738480",
  2983 => x"8080f52d",
  2984 => x"7081ff06",
  2985 => x"53535470",
  2986 => x"742ea338",
  2987 => x"7181ff06",
  2988 => x"5170752e",
  2989 => x"09810683",
  2990 => x"38725481",
  2991 => x"13708480",
  2992 => x"8080f52d",
  2993 => x"7081ff06",
  2994 => x"53535370",
  2995 => x"df387383",
  2996 => x"ffe0800c",
  2997 => x"0294050d",
  2998 => x"0402e805",
  2999 => x"0d77797b",
  3000 => x"72720783",
  3001 => x"06545456",
  3002 => x"5670802e",
  3003 => x"aa387476",
  3004 => x"5253ff12",
  3005 => x"5271ff2e",
  3006 => x"80f43872",
  3007 => x"70810554",
  3008 => x"84808080",
  3009 => x"f52d7170",
  3010 => x"81055384",
  3011 => x"808081b7",
  3012 => x"2d848080",
  3013 => x"ddf20474",
  3014 => x"7673822a",
  3015 => x"ff055354",
  3016 => x"5470ff2e",
  3017 => x"96387370",
  3018 => x"84055508",
  3019 => x"73708405",
  3020 => x"550cff11",
  3021 => x"51848080",
  3022 => x"dea10471",
  3023 => x"fc067016",
  3024 => x"55760572",
  3025 => x"8306ff05",
  3026 => x"525370ff",
  3027 => x"2ea03873",
  3028 => x"70810555",
  3029 => x"84808080",
  3030 => x"f52d7370",
  3031 => x"81055584",
  3032 => x"808081b7",
  3033 => x"2dff1151",
  3034 => x"848080de",
  3035 => x"ca047583",
  3036 => x"ffe0800c",
  3037 => x"0298050d",
  3038 => x"0402f005",
  3039 => x"0d757078",
  3040 => x"ff1b5454",
  3041 => x"545470ff",
  3042 => x"2ea03871",
  3043 => x"70810553",
  3044 => x"84808080",
  3045 => x"f52d7370",
  3046 => x"81055584",
  3047 => x"808081b7",
  3048 => x"2dff1151",
  3049 => x"848080df",
  3050 => x"86047383",
  3051 => x"ffe0800c",
  3052 => x"0290050d",
  3053 => x"0402ec05",
  3054 => x"0d787779",
  3055 => x"53545284",
  3056 => x"8080dfd3",
  3057 => x"04ff1252",
  3058 => x"71ff2e9c",
  3059 => x"38811381",
  3060 => x"12525370",
  3061 => x"84808080",
  3062 => x"f52d7384",
  3063 => x"808080f5",
  3064 => x"2d565473",
  3065 => x"752ede38",
  3066 => x"72848080",
  3067 => x"80f52d71",
  3068 => x"84808080",
  3069 => x"f52d7171",
  3070 => x"3183ffe0",
  3071 => x"800c5253",
  3072 => x"0294050d",
  3073 => x"0402f005",
  3074 => x"0d767877",
  3075 => x"54525384",
  3076 => x"8080e0a0",
  3077 => x"04ff1151",
  3078 => x"70ff2e94",
  3079 => x"38811252",
  3080 => x"71848080",
  3081 => x"80f52d54",
  3082 => x"72742e09",
  3083 => x"8106e638",
  3084 => x"71728480",
  3085 => x"8080f52d",
  3086 => x"53517272",
  3087 => x"2e833880",
  3088 => x"517083ff",
  3089 => x"e0800c02",
  3090 => x"90050d04",
  3091 => x"02f0050d",
  3092 => x"757771ff",
  3093 => x"1b545455",
  3094 => x"5370ff2e",
  3095 => x"96387372",
  3096 => x"70810554",
  3097 => x"84808081",
  3098 => x"b72dff11",
  3099 => x"51848080",
  3100 => x"e0d90472",
  3101 => x"83ffe080",
  3102 => x"0c029005",
  3103 => x"0d0402f0",
  3104 => x"050d7552",
  3105 => x"848080e1",
  3106 => x"8d048112",
  3107 => x"52807284",
  3108 => x"808080f5",
  3109 => x"2d7081ff",
  3110 => x"06535454",
  3111 => x"70742e83",
  3112 => x"38815470",
  3113 => x"a02e8438",
  3114 => x"73e03872",
  3115 => x"81ff0651",
  3116 => x"70a02e09",
  3117 => x"81069238",
  3118 => x"81127084",
  3119 => x"808080f5",
  3120 => x"2d525284",
  3121 => x"8080e1b0",
  3122 => x"04718480",
  3123 => x"8080f52d",
  3124 => x"70545170",
  3125 => x"802e8338",
  3126 => x"71537283",
  3127 => x"ffe0800c",
  3128 => x"0290050d",
  3129 => x"0402e805",
  3130 => x"0d777957",
  3131 => x"55805473",
  3132 => x"7524b338",
  3133 => x"75742953",
  3134 => x"72752e09",
  3135 => x"81068938",
  3136 => x"80538480",
  3137 => x"80e2a604",
  3138 => x"74732591",
  3139 => x"38737629",
  3140 => x"76317571",
  3141 => x"31515384",
  3142 => x"8080e2a6",
  3143 => x"04811454",
  3144 => x"848080e1",
  3145 => x"ef047283",
  3146 => x"ffe0800c",
  3147 => x"0298050d",
  3148 => x"0402e005",
  3149 => x"0d797b58",
  3150 => x"56807059",
  3151 => x"54775377",
  3152 => x"762eb638",
  3153 => x"77762499",
  3154 => x"38811477",
  3155 => x"19595475",
  3156 => x"7427ea38",
  3157 => x"72547485",
  3158 => x"249f3884",
  3159 => x"8080e2f7",
  3160 => x"04737729",
  3161 => x"77317671",
  3162 => x"31902b70",
  3163 => x"902c5156",
  3164 => x"53848080",
  3165 => x"e2d40472",
  3166 => x"547383ff",
  3167 => x"e0800c02",
  3168 => x"a0050d04",
  3169 => x"02f8050d",
  3170 => x"74527351",
  3171 => x"848080e2",
  3172 => x"b12d0288",
  3173 => x"050d0402",
  3174 => x"f8050d74",
  3175 => x"52735184",
  3176 => x"8080e1e5",
  3177 => x"2d028805",
  3178 => x"0d0402cc",
  3179 => x"050d8480",
  3180 => x"80e9e451",
  3181 => x"84808082",
  3182 => x"e32d8480",
  3183 => x"80e9f451",
  3184 => x"84808082",
  3185 => x"e32d8480",
  3186 => x"80ea8c51",
  3187 => x"84808082",
  3188 => x"e32d8480",
  3189 => x"8087be2d",
  3190 => x"83ffe080",
  3191 => x"0881ce38",
  3192 => x"8480808d",
  3193 => x"b72d8480",
  3194 => x"80b3a62d",
  3195 => x"84808090",
  3196 => x"dc528480",
  3197 => x"8090aa51",
  3198 => x"848080b3",
  3199 => x"f42d83ff",
  3200 => x"e0800880",
  3201 => x"2e80c438",
  3202 => x"848080ea",
  3203 => x"a0518480",
  3204 => x"8082e32d",
  3205 => x"81558480",
  3206 => x"80e6f904",
  3207 => x"83ffe080",
  3208 => x"08549080",
  3209 => x"80538152",
  3210 => x"80c0c084",
  3211 => x"51848080",
  3212 => x"b9c62d83",
  3213 => x"ffe08008",
  3214 => x"52848080",
  3215 => x"eabc5184",
  3216 => x"808082e3",
  3217 => x"2d848080",
  3218 => x"e5dc0484",
  3219 => x"8080ead0",
  3220 => x"51848080",
  3221 => x"82e32d84",
  3222 => x"8080eaec",
  3223 => x"51848080",
  3224 => x"c2ae2d84",
  3225 => x"8080eaf0",
  3226 => x"51848080",
  3227 => x"82e32d80",
  3228 => x"53885202",
  3229 => x"a8057052",
  3230 => x"55848080",
  3231 => x"86ae2d84",
  3232 => x"8080eb80",
  3233 => x"52745184",
  3234 => x"8080b596",
  3235 => x"2d83ffe0",
  3236 => x"80085a83",
  3237 => x"ffe08008",
  3238 => x"ff823884",
  3239 => x"8080eb84",
  3240 => x"51848080",
  3241 => x"82e32d84",
  3242 => x"8080e4e3",
  3243 => x"04848080",
  3244 => x"eba05184",
  3245 => x"808082e3",
  3246 => x"2d805388",
  3247 => x"5202a805",
  3248 => x"55745184",
  3249 => x"808086ae",
  3250 => x"2d748480",
  3251 => x"80ebcc2e",
  3252 => x"8b388053",
  3253 => x"88528480",
  3254 => x"80e5c104",
  3255 => x"80597882",
  3256 => x"2b80c0c0",
  3257 => x"87118480",
  3258 => x"8080f52d",
  3259 => x"80c0c086",
  3260 => x"12848080",
  3261 => x"80f52d71",
  3262 => x"982b7190",
  3263 => x"2b0780c0",
  3264 => x"c0851484",
  3265 => x"808080f5",
  3266 => x"2d70882b",
  3267 => x"720780c0",
  3268 => x"c0841684",
  3269 => x"808080f5",
  3270 => x"2d710770",
  3271 => x"882a83fe",
  3272 => x"80067072",
  3273 => x"982a0772",
  3274 => x"882b87fc",
  3275 => x"80800671",
  3276 => x"0773982b",
  3277 => x"07790c51",
  3278 => x"53515253",
  3279 => x"58595758",
  3280 => x"81195983",
  3281 => x"ffff7925",
  3282 => x"ff943884",
  3283 => x"8080ebd0",
  3284 => x"51848080",
  3285 => x"82e32d79",
  3286 => x"51848080",
  3287 => x"b8cf2d84",
  3288 => x"8080b4db",
  3289 => x"2d848080",
  3290 => x"80932d84",
  3291 => x"8080ebdc",
  3292 => x"51848080",
  3293 => x"82e32d80",
  3294 => x"557483ff",
  3295 => x"e0800c02",
  3296 => x"b4050d04",
  3297 => x"00ffffff",
  3298 => x"ff00ffff",
  3299 => x"ffff00ff",
  3300 => x"ffffff00",
  3301 => x"08200800",
  3302 => x"434d4438",
  3303 => x"5f342072",
  3304 => x"6573706f",
  3305 => x"6e73653a",
  3306 => x"2025640a",
  3307 => x"00000000",
  3308 => x"53444843",
  3309 => x"20496e69",
  3310 => x"7469616c",
  3311 => x"697a6174",
  3312 => x"696f6e20",
  3313 => x"6572726f",
  3314 => x"72210a00",
  3315 => x"434d4435",
  3316 => x"38202564",
  3317 => x"0a202000",
  3318 => x"52656164",
  3319 => x"20636f6d",
  3320 => x"6d616e64",
  3321 => x"20666169",
  3322 => x"6c656420",
  3323 => x"61742025",
  3324 => x"64202825",
  3325 => x"64290a00",
  3326 => x"4641545f",
  3327 => x"46533a20",
  3328 => x"4572726f",
  3329 => x"7220636f",
  3330 => x"756c6420",
  3331 => x"6e6f7420",
  3332 => x"6c6f6164",
  3333 => x"20464154",
  3334 => x"20646574",
  3335 => x"61696c73",
  3336 => x"20282564",
  3337 => x"29210d0a",
  3338 => x"00000000",
  3339 => x"2573203c",
  3340 => x"4449523e",
  3341 => x"0d0a0000",
  3342 => x"2573205b",
  3343 => x"25642062",
  3344 => x"79746573",
  3345 => x"5d0d0a00",
  3346 => x"46415420",
  3347 => x"64657461",
  3348 => x"696c733a",
  3349 => x"0d0a0000",
  3350 => x"46415433",
  3351 => x"32000000",
  3352 => x"46415431",
  3353 => x"36000000",
  3354 => x"20547970",
  3355 => x"65203d25",
  3356 => x"73000000",
  3357 => x"20526f6f",
  3358 => x"74204469",
  3359 => x"72204669",
  3360 => x"72737420",
  3361 => x"436c7573",
  3362 => x"74657220",
  3363 => x"3d202578",
  3364 => x"0d0a0000",
  3365 => x"20464154",
  3366 => x"20426567",
  3367 => x"696e204c",
  3368 => x"4241203d",
  3369 => x"20307825",
  3370 => x"780d0a00",
  3371 => x"20436c75",
  3372 => x"73746572",
  3373 => x"20426567",
  3374 => x"696e204c",
  3375 => x"4241203d",
  3376 => x"20307825",
  3377 => x"780d0a00",
  3378 => x"20536563",
  3379 => x"746f7273",
  3380 => x"20506572",
  3381 => x"20436c75",
  3382 => x"73746572",
  3383 => x"203d2025",
  3384 => x"640d0a00",
  3385 => x"426f6f74",
  3386 => x"206f7074",
  3387 => x"696f6e73",
  3388 => x"3a0a0000",
  3389 => x"30203a20",
  3390 => x"426f6f74",
  3391 => x"2066726f",
  3392 => x"6d205344",
  3393 => x"20636172",
  3394 => x"640a0000",
  3395 => x"31203a20",
  3396 => x"426f6f74",
  3397 => x"2066726f",
  3398 => x"6d204a54",
  3399 => x"41470a00",
  3400 => x"4552524f",
  3401 => x"523a204d",
  3402 => x"65646961",
  3403 => x"20617474",
  3404 => x"61636820",
  3405 => x"6661696c",
  3406 => x"65640a00",
  3407 => x"0a202564",
  3408 => x"20627974",
  3409 => x"65732072",
  3410 => x"6561640a",
  3411 => x"00000000",
  3412 => x"4c697374",
  3413 => x"696e6720",
  3414 => x"64697265",
  3415 => x"63746f72",
  3416 => x"6965732e",
  3417 => x"2e2e0a0a",
  3418 => x"00000000",
  3419 => x"2f000000",
  3420 => x"0a415050",
  3421 => x"2046494c",
  3422 => x"45203e3e",
  3423 => x"20000000",
  3424 => x"72620000",
  3425 => x"4552524f",
  3426 => x"523a2052",
  3427 => x"65616420",
  3428 => x"66696c65",
  3429 => x"20666169",
  3430 => x"6c65640a",
  3431 => x"00000000",
  3432 => x"426f6f74",
  3433 => x"696e6720",
  3434 => x"66726f6d",
  3435 => x"204a5441",
  3436 => x"472c2077",
  3437 => x"61697469",
  3438 => x"6e672066",
  3439 => x"6f722075",
  3440 => x"706c6f61",
  3441 => x"6465720a",
  3442 => x"00000000",
  3443 => x"454e4400",
  3444 => x"0a0a456e",
  3445 => x"642e2e2e",
  3446 => x"200a0000",
  3447 => x"73687574",
  3448 => x"646f776e",
  3449 => x"2e0a0000",
others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;

		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end rtl;

