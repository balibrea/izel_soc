--
-- (C) 2018, ZPUROMGEN, Yosel de Jesus Balibrea Lastre.
--           Automatically Generated ROM file
--           Please do NOT CHANGE!
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity prog_mem is
generic
(
maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
);
port (
		clk : in std_logic;
		areset : in std_logic := '0';
		from_zpu : in ZPU_ToROM;
		to_zpu : out ZPU_FromROM
		);
end prog_mem;

architecture rtl of prog_mem is

	type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

	shared variable ram : ram_type := (
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080e7c8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff2",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"8080e3d6",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c32d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870892a",
   171 => x"70810651",
   172 => x"515170f3",
   173 => x"3871c00c",
   174 => x"7183ffe0",
   175 => x"800c0288",
   176 => x"050d0402",
   177 => x"e8050d80",
   178 => x"78575575",
   179 => x"70840557",
   180 => x"08538054",
   181 => x"72982a73",
   182 => x"882b5452",
   183 => x"71802ea0",
   184 => x"38c00870",
   185 => x"892a7081",
   186 => x"06515151",
   187 => x"70f33871",
   188 => x"c00c8115",
   189 => x"81155555",
   190 => x"837425d8",
   191 => x"3871cc38",
   192 => x"7483ffe0",
   193 => x"800c0298",
   194 => x"050d0402",
   195 => x"fc050dc0",
   196 => x"0870882a",
   197 => x"70810651",
   198 => x"515170f3",
   199 => x"38c00870",
   200 => x"81ff0683",
   201 => x"ffe0800c",
   202 => x"51028405",
   203 => x"0d0402e4",
   204 => x"050d787a",
   205 => x"7c585855",
   206 => x"80547377",
   207 => x"2580f438",
   208 => x"84808086",
   209 => x"8b2d83ff",
   210 => x"e0800881",
   211 => x"ff065372",
   212 => x"882e0981",
   213 => x"06a33880",
   214 => x"7425df38",
   215 => x"75802e8d",
   216 => x"38848080",
   217 => x"e7d85184",
   218 => x"808085c3",
   219 => x"2dff15ff",
   220 => x"15555584",
   221 => x"808086ba",
   222 => x"04728d2e",
   223 => x"b638e013",
   224 => x"527180de",
   225 => x"26ffb338",
   226 => x"75802e92",
   227 => x"38c00870",
   228 => x"892a7081",
   229 => x"06515152",
   230 => x"71f33872",
   231 => x"c00c7275",
   232 => x"70810557",
   233 => x"84808081",
   234 => x"b72d8114",
   235 => x"54848080",
   236 => x"86ba0480",
   237 => x"75848080",
   238 => x"81b72d73",
   239 => x"83ffe080",
   240 => x"0c029c05",
   241 => x"0d0402d0",
   242 => x"050d8070",
   243 => x"57578177",
   244 => x"54588852",
   245 => x"02a40570",
   246 => x"52598480",
   247 => x"8086ae2d",
   248 => x"76557419",
   249 => x"70848080",
   250 => x"80f52d89",
   251 => x"0bd01227",
   252 => x"78058118",
   253 => x"58585154",
   254 => x"877525e6",
   255 => x"38807625",
   256 => x"a63802a3",
   257 => x"05557515",
   258 => x"70848080",
   259 => x"80f52dd0",
   260 => x"117a2979",
   261 => x"057a8829",
   262 => x"7b1005ff",
   263 => x"1a5a5b59",
   264 => x"51547580",
   265 => x"24e03876",
   266 => x"83ffe080",
   267 => x"0c02b005",
   268 => x"0d0402f4",
   269 => x"050dd452",
   270 => x"81ff720c",
   271 => x"71085381",
   272 => x"ff720c72",
   273 => x"882b83fe",
   274 => x"80067208",
   275 => x"7081ff06",
   276 => x"51525381",
   277 => x"ff720c72",
   278 => x"7107882b",
   279 => x"72087081",
   280 => x"ff065152",
   281 => x"5381ff72",
   282 => x"0c727107",
   283 => x"882b7208",
   284 => x"7081ff06",
   285 => x"720783ff",
   286 => x"e0800c52",
   287 => x"53028c05",
   288 => x"0d0402f4",
   289 => x"050d7476",
   290 => x"7181ff06",
   291 => x"d40c5353",
   292 => x"83fff2e4",
   293 => x"08853871",
   294 => x"892b5271",
   295 => x"982ad40c",
   296 => x"71902a70",
   297 => x"81ff06d4",
   298 => x"0c517188",
   299 => x"2a7081ff",
   300 => x"06d40c51",
   301 => x"7181ff06",
   302 => x"d40c7290",
   303 => x"2a7081ff",
   304 => x"06d40c51",
   305 => x"d4087081",
   306 => x"ff065151",
   307 => x"82b8bf52",
   308 => x"7081ff2e",
   309 => x"09810694",
   310 => x"3881ff0b",
   311 => x"d40cd408",
   312 => x"7081ff06",
   313 => x"ff145451",
   314 => x"5171e538",
   315 => x"7083ffe0",
   316 => x"800c028c",
   317 => x"050d0402",
   318 => x"fc050d81",
   319 => x"c75181ff",
   320 => x"0bd40cff",
   321 => x"11517080",
   322 => x"25f43802",
   323 => x"84050d04",
   324 => x"02f0050d",
   325 => x"84808089",
   326 => x"f72d819c",
   327 => x"9f538052",
   328 => x"87fc80f7",
   329 => x"51848080",
   330 => x"89822d83",
   331 => x"ffe08008",
   332 => x"5483ffe0",
   333 => x"8008812e",
   334 => x"098106ae",
   335 => x"3881ff0b",
   336 => x"d40c820a",
   337 => x"52849c80",
   338 => x"e9518480",
   339 => x"8089822d",
   340 => x"83ffe080",
   341 => x"088e3881",
   342 => x"ff0bd40c",
   343 => x"73538480",
   344 => x"808af104",
   345 => x"84808089",
   346 => x"f72dff13",
   347 => x"5372ffae",
   348 => x"387283ff",
   349 => x"e0800c02",
   350 => x"90050d04",
   351 => x"02f4050d",
   352 => x"81ff0bd4",
   353 => x"0c935380",
   354 => x"5287fc80",
   355 => x"c1518480",
   356 => x"8089822d",
   357 => x"83ffe080",
   358 => x"088e3881",
   359 => x"ff0bd40c",
   360 => x"81538480",
   361 => x"808bb404",
   362 => x"84808089",
   363 => x"f72dff13",
   364 => x"5372d438",
   365 => x"7283ffe0",
   366 => x"800c028c",
   367 => x"050d0402",
   368 => x"f0050d84",
   369 => x"808089f7",
   370 => x"2d83aa52",
   371 => x"849c80c8",
   372 => x"51848080",
   373 => x"89822d83",
   374 => x"ffe08008",
   375 => x"812e0981",
   376 => x"06a93884",
   377 => x"808088b2",
   378 => x"2d83ffe0",
   379 => x"800883ff",
   380 => x"ff065372",
   381 => x"83aa2ebb",
   382 => x"3883ffe0",
   383 => x"80085284",
   384 => x"8080e7dc",
   385 => x"51848080",
   386 => x"82e32d84",
   387 => x"80808afc",
   388 => x"2d848080",
   389 => x"8cab0481",
   390 => x"54848080",
   391 => x"8db40484",
   392 => x"8080e7f4",
   393 => x"51848080",
   394 => x"82e32d80",
   395 => x"54848080",
   396 => x"8db40481",
   397 => x"ff0bd40c",
   398 => x"b1538480",
   399 => x"808a902d",
   400 => x"83ffe080",
   401 => x"08802e80",
   402 => x"dc388052",
   403 => x"87fc80fa",
   404 => x"51848080",
   405 => x"89822d83",
   406 => x"ffe08008",
   407 => x"b63881ff",
   408 => x"0bd40cd4",
   409 => x"085381ff",
   410 => x"0bd40c81",
   411 => x"ff0bd40c",
   412 => x"81ff0bd4",
   413 => x"0c81ff0b",
   414 => x"d40c7286",
   415 => x"2a708106",
   416 => x"83ffe080",
   417 => x"08565153",
   418 => x"72802ea8",
   419 => x"38848080",
   420 => x"8c970483",
   421 => x"ffe08008",
   422 => x"52848080",
   423 => x"e8905184",
   424 => x"808082e3",
   425 => x"2d72822e",
   426 => x"fef538ff",
   427 => x"135372ff",
   428 => x"89387254",
   429 => x"7383ffe0",
   430 => x"800c0290",
   431 => x"050d0402",
   432 => x"f4050d81",
   433 => x"0b83fff2",
   434 => x"e40cd008",
   435 => x"708f2a70",
   436 => x"81065151",
   437 => x"5372f338",
   438 => x"72d00c84",
   439 => x"808089f7",
   440 => x"2dd00870",
   441 => x"8f2a7081",
   442 => x"06515153",
   443 => x"72f33881",
   444 => x"0bd00c87",
   445 => x"53805284",
   446 => x"d480c051",
   447 => x"84808089",
   448 => x"822d83ff",
   449 => x"e0800881",
   450 => x"2e973872",
   451 => x"822e0981",
   452 => x"06893880",
   453 => x"53848080",
   454 => x"8ee204ff",
   455 => x"135372d5",
   456 => x"38848080",
   457 => x"8bbf2d83",
   458 => x"ffe08008",
   459 => x"83fff2e4",
   460 => x"0c83ffe0",
   461 => x"80088e38",
   462 => x"815287fc",
   463 => x"80d05184",
   464 => x"80808982",
   465 => x"2d81ff0b",
   466 => x"d40cd008",
   467 => x"708f2a70",
   468 => x"81065151",
   469 => x"5372f338",
   470 => x"72d00c81",
   471 => x"ff0bd40c",
   472 => x"81537283",
   473 => x"ffe0800c",
   474 => x"028c050d",
   475 => x"04800b83",
   476 => x"ffe0800c",
   477 => x"0402e005",
   478 => x"0d797b57",
   479 => x"57805881",
   480 => x"ff0bd40c",
   481 => x"d008708f",
   482 => x"2a708106",
   483 => x"51515473",
   484 => x"f3388281",
   485 => x"0bd00c81",
   486 => x"ff0bd40c",
   487 => x"765287fc",
   488 => x"80d15184",
   489 => x"80808982",
   490 => x"2d80dbc6",
   491 => x"df5583ff",
   492 => x"e0800880",
   493 => x"2e9b3883",
   494 => x"ffe08008",
   495 => x"53765284",
   496 => x"8080e89c",
   497 => x"51848080",
   498 => x"82e32d84",
   499 => x"808090a7",
   500 => x"0481ff0b",
   501 => x"d40cd408",
   502 => x"7081ff06",
   503 => x"51547381",
   504 => x"fe2e0981",
   505 => x"06a53880",
   506 => x"ff548480",
   507 => x"8088b22d",
   508 => x"83ffe080",
   509 => x"08767084",
   510 => x"05580cff",
   511 => x"14547380",
   512 => x"25e83881",
   513 => x"58848080",
   514 => x"909104ff",
   515 => x"155574c1",
   516 => x"3881ff0b",
   517 => x"d40cd008",
   518 => x"708f2a70",
   519 => x"81065151",
   520 => x"5473f338",
   521 => x"73d00c77",
   522 => x"83ffe080",
   523 => x"0c02a005",
   524 => x"0d0402ec",
   525 => x"050d7678",
   526 => x"7a555555",
   527 => x"80732798",
   528 => x"38735274",
   529 => x"51848080",
   530 => x"8ef52d81",
   531 => x"15848015",
   532 => x"ff155555",
   533 => x"5572ea38",
   534 => x"810b83ff",
   535 => x"e0800c02",
   536 => x"94050d04",
   537 => x"02fc050d",
   538 => x"74518071",
   539 => x"278738ff",
   540 => x"115170fb",
   541 => x"38810b83",
   542 => x"ffe0800c",
   543 => x"0284050d",
   544 => x"0402fc05",
   545 => x"0d7270ff",
   546 => x"b40c83ff",
   547 => x"e0800c02",
   548 => x"84050d04",
   549 => x"ffb40883",
   550 => x"ffe0800c",
   551 => x"04c80883",
   552 => x"ffe0800c",
   553 => x"0402ec05",
   554 => x"0d765480",
   555 => x"0b84d415",
   556 => x"0cff0b88",
   557 => x"d8150c80",
   558 => x"0b88dc15",
   559 => x"0c84d814",
   560 => x"55848053",
   561 => x"80527451",
   562 => x"848080e0",
   563 => x"f82d800b",
   564 => x"88e0150c",
   565 => x"84d41408",
   566 => x"88e4150c",
   567 => x"7484d415",
   568 => x"0c029405",
   569 => x"0d0402d8",
   570 => x"050d7b7d",
   571 => x"70565855",
   572 => x"76802e80",
   573 => x"d0388484",
   574 => x"1708802e",
   575 => x"80c538b8",
   576 => x"15085978",
   577 => x"802eb638",
   578 => x"810b8480",
   579 => x"18087094",
   580 => x"18083172",
   581 => x"11a01908",
   582 => x"59575859",
   583 => x"5a747427",
   584 => x"85387476",
   585 => x"315a7953",
   586 => x"76527751",
   587 => x"782d83ff",
   588 => x"e0800854",
   589 => x"83ffe080",
   590 => x"08802e89",
   591 => x"38800b84",
   592 => x"84180c81",
   593 => x"547383ff",
   594 => x"e0800c02",
   595 => x"a8050d04",
   596 => x"02e0050d",
   597 => x"797b5957",
   598 => x"800b84d4",
   599 => x"18085656",
   600 => x"74762e80",
   601 => x"db388480",
   602 => x"15085473",
   603 => x"78268938",
   604 => x"81145473",
   605 => x"7826ae38",
   606 => x"848c1508",
   607 => x"54739638",
   608 => x"75802e8c",
   609 => x"3873848c",
   610 => x"170c8480",
   611 => x"80939504",
   612 => x"7584d418",
   613 => x"0c74848c",
   614 => x"16085656",
   615 => x"74c83884",
   616 => x"808093c0",
   617 => x"0474802e",
   618 => x"97387784",
   619 => x"80160831",
   620 => x"892b7505",
   621 => x"8488160c",
   622 => x"74548480",
   623 => x"8094a204",
   624 => x"84d41708",
   625 => x"848c170c",
   626 => x"7584d418",
   627 => x"0c848416",
   628 => x"08802e9a",
   629 => x"38755276",
   630 => x"51848080",
   631 => x"91e62d83",
   632 => x"ffe08008",
   633 => x"5483ffe0",
   634 => x"8008802e",
   635 => x"b5387784",
   636 => x"80170c81",
   637 => x"53755284",
   638 => x"80160851",
   639 => x"b4170854",
   640 => x"732d83ff",
   641 => x"e0800893",
   642 => x"38ff0b84",
   643 => x"80170c83",
   644 => x"ffe08008",
   645 => x"54848080",
   646 => x"94a20475",
   647 => x"8488170c",
   648 => x"75547383",
   649 => x"ffe0800c",
   650 => x"02a0050d",
   651 => x"0402f005",
   652 => x"0d7584d4",
   653 => x"11085454",
   654 => x"72802eb1",
   655 => x"38848413",
   656 => x"08802e9e",
   657 => x"38725273",
   658 => x"51848080",
   659 => x"91e62d83",
   660 => x"ffe08008",
   661 => x"8d3883ff",
   662 => x"e0800853",
   663 => x"84808094",
   664 => x"ef04848c",
   665 => x"13085384",
   666 => x"808094b8",
   667 => x"04815372",
   668 => x"83ffe080",
   669 => x"0c029005",
   670 => x"0d0402e8",
   671 => x"050d7779",
   672 => x"55567383",
   673 => x"38825473",
   674 => x"882a53b0",
   675 => x"1608802e",
   676 => x"85387387",
   677 => x"2a539416",
   678 => x"08135275",
   679 => x"51848080",
   680 => x"92d02dff",
   681 => x"5583ffe0",
   682 => x"8008802e",
   683 => x"819a3883",
   684 => x"ffe08008",
   685 => x"84880508",
   686 => x"55b01608",
   687 => x"b2387288",
   688 => x"2b747131",
   689 => x"107083ff",
   690 => x"fe061781",
   691 => x"11848080",
   692 => x"80f52d71",
   693 => x"84808080",
   694 => x"f52d7182",
   695 => x"802905fc",
   696 => x"80881153",
   697 => x"58585151",
   698 => x"53848080",
   699 => x"96bf0472",
   700 => x"872b7471",
   701 => x"31822b83",
   702 => x"fffc0616",
   703 => x"83118480",
   704 => x"8080f52d",
   705 => x"82128480",
   706 => x"8080f52d",
   707 => x"7181800a",
   708 => x"29718480",
   709 => x"80290581",
   710 => x"14848080",
   711 => x"80f52d70",
   712 => x"82802912",
   713 => x"75848080",
   714 => x"80f52d56",
   715 => x"7505f00a",
   716 => x"06ff8080",
   717 => x"80881153",
   718 => x"55535459",
   719 => x"575553ff",
   720 => x"55877327",
   721 => x"83387355",
   722 => x"7483ffe0",
   723 => x"800c0298",
   724 => x"050d0402",
   725 => x"e0050d79",
   726 => x"7b5856b0",
   727 => x"1608802e",
   728 => x"81ba3898",
   729 => x"16848080",
   730 => x"80e02d9c",
   731 => x"17080552",
   732 => x"75518480",
   733 => x"8092d02d",
   734 => x"83ffe080",
   735 => x"085883ff",
   736 => x"e0800880",
   737 => x"2e819538",
   738 => x"83ffe080",
   739 => x"08848805",
   740 => x"08547683",
   741 => x"ec158480",
   742 => x"8081b72d",
   743 => x"83ffe080",
   744 => x"08848805",
   745 => x"0877882a",
   746 => x"55557383",
   747 => x"ed168480",
   748 => x"8081b72d",
   749 => x"83ffe080",
   750 => x"08848805",
   751 => x"0877902a",
   752 => x"55557383",
   753 => x"ee168480",
   754 => x"8081b72d",
   755 => x"83ffe080",
   756 => x"08848805",
   757 => x"0877982a",
   758 => x"55557383",
   759 => x"ef168480",
   760 => x"8081b72d",
   761 => x"810b83ff",
   762 => x"e0800884",
   763 => x"84050c76",
   764 => x"a4170cb8",
   765 => x"16085473",
   766 => x"802e9538",
   767 => x"815383ff",
   768 => x"e0800852",
   769 => x"83ffe080",
   770 => x"08848005",
   771 => x"0851732d",
   772 => x"ff0b8480",
   773 => x"190c800b",
   774 => x"8484190c",
   775 => x"02a0050d",
   776 => x"0402d005",
   777 => x"0d7d5780",
   778 => x"705956a0",
   779 => x"1708762e",
   780 => x"81ba3894",
   781 => x"17081852",
   782 => x"76518480",
   783 => x"8092d02d",
   784 => x"83ffe080",
   785 => x"08802e81",
   786 => x"a338800b",
   787 => x"b0180883",
   788 => x"ffe08008",
   789 => x"84880508",
   790 => x"5b5b5574",
   791 => x"83ffff06",
   792 => x"5379ad38",
   793 => x"72198111",
   794 => x"84808080",
   795 => x"f52d7184",
   796 => x"808080f5",
   797 => x"2d718280",
   798 => x"29057081",
   799 => x"05097080",
   800 => x"251a821a",
   801 => x"5a5a5152",
   802 => x"55538480",
   803 => x"8099da04",
   804 => x"72198311",
   805 => x"84808080",
   806 => x"f52d8212",
   807 => x"84808080",
   808 => x"f52d7181",
   809 => x"800a2971",
   810 => x"84808029",
   811 => x"05811484",
   812 => x"808080f5",
   813 => x"2d708280",
   814 => x"29127584",
   815 => x"808080f5",
   816 => x"2d710570",
   817 => x"81050970",
   818 => x"72078025",
   819 => x"7e05841e",
   820 => x"5e5e5751",
   821 => x"5253575d",
   822 => x"5d5383ff",
   823 => x"7527fefb",
   824 => x"38811858",
   825 => x"a0170878",
   826 => x"26fec838",
   827 => x"7583ffe0",
   828 => x"800c02b0",
   829 => x"050d0402",
   830 => x"ec050d76",
   831 => x"538054ff",
   832 => x"5272742e",
   833 => x"81963872",
   834 => x"84808080",
   835 => x"f52d5170",
   836 => x"af2e0981",
   837 => x"068c3870",
   838 => x"81145455",
   839 => x"8480809a",
   840 => x"cc048113",
   841 => x"84808080",
   842 => x"f52d5170",
   843 => x"ba2e9638",
   844 => x"82138480",
   845 => x"8080f52d",
   846 => x"51ff5270",
   847 => x"80dc2e09",
   848 => x"810680d8",
   849 => x"3880dc0b",
   850 => x"83145455",
   851 => x"72848080",
   852 => x"80f52d70",
   853 => x"81ff0652",
   854 => x"5270802e",
   855 => x"bc387181",
   856 => x"ff065170",
   857 => x"802ea938",
   858 => x"7181ff06",
   859 => x"81145351",
   860 => x"70752e09",
   861 => x"81068938",
   862 => x"71538480",
   863 => x"809b9004",
   864 => x"71728480",
   865 => x"8080f52d",
   866 => x"53538480",
   867 => x"809ade04",
   868 => x"81145484",
   869 => x"80809acc",
   870 => x"04ff1452",
   871 => x"7183ffe0",
   872 => x"800c0294",
   873 => x"050d0402",
   874 => x"d0050d7d",
   875 => x"7f616358",
   876 => x"5d5d5380",
   877 => x"70748105",
   878 => x"09707607",
   879 => x"73257074",
   880 => x"7a250751",
   881 => x"51545b58",
   882 => x"ff547178",
   883 => x"2e098106",
   884 => x"81d63872",
   885 => x"84808080",
   886 => x"f52d5271",
   887 => x"af2e0981",
   888 => x"068c3871",
   889 => x"81145457",
   890 => x"8480809c",
   891 => x"98048113",
   892 => x"84808080",
   893 => x"f52d5271",
   894 => x"ba2e9638",
   895 => x"82138480",
   896 => x"8080f52d",
   897 => x"52ff5471",
   898 => x"80dc2e09",
   899 => x"81068198",
   900 => x"3880dc0b",
   901 => x"83145457",
   902 => x"72518480",
   903 => x"80d8fa2d",
   904 => x"800b83ff",
   905 => x"e0800825",
   906 => x"80cf38ff",
   907 => x"1583ffe0",
   908 => x"80085559",
   909 => x"72848080",
   910 => x"80f52d70",
   911 => x"81ff0670",
   912 => x"79327081",
   913 => x"05097080",
   914 => x"251e5e51",
   915 => x"54565679",
   916 => x"7c2e0981",
   917 => x"06993874",
   918 => x"772e9438",
   919 => x"7779258f",
   920 => x"387a1852",
   921 => x"75728480",
   922 => x"8081b72d",
   923 => x"81185881",
   924 => x"13ff1555",
   925 => x"5373ffbc",
   926 => x"387a8480",
   927 => x"8080f52d",
   928 => x"5271802e",
   929 => x"95388480",
   930 => x"80ebcc51",
   931 => x"84808085",
   932 => x"c32d8054",
   933 => x"8480809d",
   934 => x"a8048480",
   935 => x"80ebcc51",
   936 => x"84808085",
   937 => x"c32dff54",
   938 => x"7383ffe0",
   939 => x"800c02b0",
   940 => x"050d0402",
   941 => x"d8050d7b",
   942 => x"7d7f6173",
   943 => x"555c5c59",
   944 => x"57848080",
   945 => x"99f72d83",
   946 => x"ffe08008",
   947 => x"83ffe080",
   948 => x"08565683",
   949 => x"ffe08008",
   950 => x"ff2e80f2",
   951 => x"387f5478",
   952 => x"5383ffe0",
   953 => x"80085276",
   954 => x"51848080",
   955 => x"9ba72dff",
   956 => x"5583ffe0",
   957 => x"800880d6",
   958 => x"38759338",
   959 => x"83ffe080",
   960 => x"08788480",
   961 => x"8081b72d",
   962 => x"8480809e",
   963 => x"cc047651",
   964 => x"848080d8",
   965 => x"fa2d83ff",
   966 => x"e0800879",
   967 => x"52558480",
   968 => x"80d8fa2d",
   969 => x"7483ffe0",
   970 => x"80083155",
   971 => x"79752583",
   972 => x"38795574",
   973 => x"53765277",
   974 => x"51848080",
   975 => x"de852d74",
   976 => x"18ff0555",
   977 => x"80758480",
   978 => x"8081b72d",
   979 => x"80557483",
   980 => x"ffe0800c",
   981 => x"02a8050d",
   982 => x"0402e005",
   983 => x"0d797bff",
   984 => x"1e565657",
   985 => x"73ff2e80",
   986 => x"d7387684",
   987 => x"808080f5",
   988 => x"2d707684",
   989 => x"808080f5",
   990 => x"2d70ffbf",
   991 => x"14555954",
   992 => x"59537099",
   993 => x"268938a0",
   994 => x"137081ff",
   995 => x"065951ff",
   996 => x"bf125170",
   997 => x"99268938",
   998 => x"a0127081",
   999 => x"ff065751",
  1000 => x"77763151",
  1001 => x"709c3872",
  1002 => x"802e9538",
  1003 => x"71802e90",
  1004 => x"38811781",
  1005 => x"16ff1656",
  1006 => x"56578480",
  1007 => x"809ee404",
  1008 => x"80517083",
  1009 => x"ffe0800c",
  1010 => x"02a0050d",
  1011 => x"0402ec05",
  1012 => x"0d7654ff",
  1013 => x"74545572",
  1014 => x"84808080",
  1015 => x"f52d7081",
  1016 => x"ff065252",
  1017 => x"70802e9b",
  1018 => x"387181ff",
  1019 => x"065170ae",
  1020 => x"2e098106",
  1021 => x"85387274",
  1022 => x"31558113",
  1023 => x"53848080",
  1024 => x"9fd70474",
  1025 => x"83ffe080",
  1026 => x"0c029405",
  1027 => x"0d0402ec",
  1028 => x"050d7678",
  1029 => x"707113ff",
  1030 => x"05555555",
  1031 => x"5573802e",
  1032 => x"9e387184",
  1033 => x"808080f5",
  1034 => x"2d5170a0",
  1035 => x"2e098106",
  1036 => x"8e387175",
  1037 => x"31ff13ff",
  1038 => x"16565353",
  1039 => x"73e43872",
  1040 => x"83ffe080",
  1041 => x"0c029405",
  1042 => x"0d0402d4",
  1043 => x"050d7c7e",
  1044 => x"59598079",
  1045 => x"52578480",
  1046 => x"809fcd2d",
  1047 => x"83ffe080",
  1048 => x"08785256",
  1049 => x"8480809f",
  1050 => x"cd2d83ff",
  1051 => x"e0800876",
  1052 => x"09708105",
  1053 => x"09707207",
  1054 => x"7a255156",
  1055 => x"565a83ff",
  1056 => x"e08008ff",
  1057 => x"2e8c3876",
  1058 => x"5b73772e",
  1059 => x"09810681",
  1060 => x"f73883ff",
  1061 => x"e0800809",
  1062 => x"70810509",
  1063 => x"70720780",
  1064 => x"25515555",
  1065 => x"75ff2e80",
  1066 => x"e238805b",
  1067 => x"737b2e09",
  1068 => x"810681d4",
  1069 => x"3875ff2e",
  1070 => x"80d13875",
  1071 => x"19810583",
  1072 => x"ffe08008",
  1073 => x"19810571",
  1074 => x"53565784",
  1075 => x"8080d8fa",
  1076 => x"2d83ffe0",
  1077 => x"80087552",
  1078 => x"54848080",
  1079 => x"d8fa2d73",
  1080 => x"83ffe080",
  1081 => x"082e0981",
  1082 => x"06819d38",
  1083 => x"73537452",
  1084 => x"76518480",
  1085 => x"809ed92d",
  1086 => x"757a5555",
  1087 => x"83ffe080",
  1088 => x"087b2ea3",
  1089 => x"38848080",
  1090 => x"a3880478",
  1091 => x"51848080",
  1092 => x"d8fa2d83",
  1093 => x"ffe08008",
  1094 => x"78525584",
  1095 => x"8080d8fa",
  1096 => x"2d83ffe0",
  1097 => x"80085474",
  1098 => x"52785184",
  1099 => x"8080a08e",
  1100 => x"2d83ffe0",
  1101 => x"80087453",
  1102 => x"78525584",
  1103 => x"8080a08e",
  1104 => x"2d805b74",
  1105 => x"83ffe080",
  1106 => x"082e0981",
  1107 => x"06ba3883",
  1108 => x"ffe08008",
  1109 => x"53775278",
  1110 => x"51848080",
  1111 => x"9ed92d83",
  1112 => x"ffe08008",
  1113 => x"7b2e9338",
  1114 => x"848080eb",
  1115 => x"cc518480",
  1116 => x"8085c32d",
  1117 => x"848080a3",
  1118 => x"88048480",
  1119 => x"80ebcc51",
  1120 => x"84808085",
  1121 => x"c32d815b",
  1122 => x"7a83ffe0",
  1123 => x"800c02ac",
  1124 => x"050d0402",
  1125 => x"f0050d75",
  1126 => x"5372802e",
  1127 => x"80d73872",
  1128 => x"84808080",
  1129 => x"f52d7081",
  1130 => x"ff065252",
  1131 => x"70802e80",
  1132 => x"c4388113",
  1133 => x"84808080",
  1134 => x"f52d5170",
  1135 => x"af387072",
  1136 => x"81ff0652",
  1137 => x"547080dc",
  1138 => x"2e098106",
  1139 => x"83388154",
  1140 => x"70af3270",
  1141 => x"81050970",
  1142 => x"80257607",
  1143 => x"51515170",
  1144 => x"802e8938",
  1145 => x"81518480",
  1146 => x"80a3f704",
  1147 => x"81135384",
  1148 => x"8080a39f",
  1149 => x"04805170",
  1150 => x"83ffe080",
  1151 => x"0c029005",
  1152 => x"0d0402e8",
  1153 => x"050d7779",
  1154 => x"55558056",
  1155 => x"848080a4",
  1156 => x"bc047181",
  1157 => x"15555371",
  1158 => x"a02ea138",
  1159 => x"ffbf1251",
  1160 => x"70992689",
  1161 => x"38a01270",
  1162 => x"81ff0654",
  1163 => x"51727570",
  1164 => x"81055784",
  1165 => x"808081b7",
  1166 => x"2d811656",
  1167 => x"80748480",
  1168 => x"8080f52d",
  1169 => x"53517171",
  1170 => x"2e833881",
  1171 => x"51758b24",
  1172 => x"853870ff",
  1173 => x"bd388075",
  1174 => x"84808081",
  1175 => x"b72d810b",
  1176 => x"83ffe080",
  1177 => x"0c029805",
  1178 => x"0d0402e0",
  1179 => x"050d797b",
  1180 => x"7d575754",
  1181 => x"80745258",
  1182 => x"8480809f",
  1183 => x"cd2d83ff",
  1184 => x"e0800878",
  1185 => x"24527578",
  1186 => x"2e80eb38",
  1187 => x"71782e80",
  1188 => x"e5387478",
  1189 => x"2e80df38",
  1190 => x"83ffe080",
  1191 => x"08148105",
  1192 => x"70848080",
  1193 => x"80f52d54",
  1194 => x"5472782e",
  1195 => x"b938ff15",
  1196 => x"57777725",
  1197 => x"b1387281",
  1198 => x"15ffbf15",
  1199 => x"54555571",
  1200 => x"99268938",
  1201 => x"a0137081",
  1202 => x"ff065652",
  1203 => x"74767081",
  1204 => x"05588480",
  1205 => x"8081b72d",
  1206 => x"81187484",
  1207 => x"808080f5",
  1208 => x"2d545872",
  1209 => x"cc388076",
  1210 => x"84808081",
  1211 => x"b72d8152",
  1212 => x"848080a5",
  1213 => x"f8048052",
  1214 => x"7183ffe0",
  1215 => x"800c02a0",
  1216 => x"050d0402",
  1217 => x"dc050d7a",
  1218 => x"7c7e605b",
  1219 => x"55575280",
  1220 => x"705855af",
  1221 => x"72810509",
  1222 => x"7074079f",
  1223 => x"2a515259",
  1224 => x"75752e81",
  1225 => x"d9388170",
  1226 => x"72065254",
  1227 => x"70752e81",
  1228 => x"cd387281",
  1229 => x"05097074",
  1230 => x"079f2a51",
  1231 => x"51747825",
  1232 => x"81bc3870",
  1233 => x"74065170",
  1234 => x"752e81b2",
  1235 => x"38718480",
  1236 => x"8080f52d",
  1237 => x"5170752e",
  1238 => x"b338fe18",
  1239 => x"54747425",
  1240 => x"ab387081",
  1241 => x"13535770",
  1242 => x"80dc2e09",
  1243 => x"81068338",
  1244 => x"70597673",
  1245 => x"70810555",
  1246 => x"84808081",
  1247 => x"b72d8115",
  1248 => x"72848080",
  1249 => x"80f52d52",
  1250 => x"5570d238",
  1251 => x"7680dc32",
  1252 => x"70810509",
  1253 => x"7072079f",
  1254 => x"2a515252",
  1255 => x"76af2e92",
  1256 => x"3870802e",
  1257 => x"8d387873",
  1258 => x"70810555",
  1259 => x"84808081",
  1260 => x"b72d7584",
  1261 => x"808080f5",
  1262 => x"2d7081ff",
  1263 => x"06525270",
  1264 => x"802eab38",
  1265 => x"ff185474",
  1266 => x"7425a338",
  1267 => x"81165671",
  1268 => x"73708105",
  1269 => x"55848080",
  1270 => x"81b72d81",
  1271 => x"15768480",
  1272 => x"8080f52d",
  1273 => x"7081ff06",
  1274 => x"53535570",
  1275 => x"da388073",
  1276 => x"84808081",
  1277 => x"b72d8151",
  1278 => x"848080a8",
  1279 => x"80048051",
  1280 => x"7083ffe0",
  1281 => x"800c02a4",
  1282 => x"050d0402",
  1283 => x"fc050d72",
  1284 => x"51807184",
  1285 => x"808081b7",
  1286 => x"2d028405",
  1287 => x"0d0402fc",
  1288 => x"050d728b",
  1289 => x"11848080",
  1290 => x"80f52d70",
  1291 => x"8f06708f",
  1292 => x"32708105",
  1293 => x"09708025",
  1294 => x"83ffe080",
  1295 => x"0c515151",
  1296 => x"51510284",
  1297 => x"050d0402",
  1298 => x"f8050d73",
  1299 => x"8b118480",
  1300 => x"8080f52d",
  1301 => x"5252708f",
  1302 => x"2ea43871",
  1303 => x"84808080",
  1304 => x"f52d5271",
  1305 => x"802e9738",
  1306 => x"7181e52e",
  1307 => x"91387088",
  1308 => x"2e8c3870",
  1309 => x"86065181",
  1310 => x"5270802e",
  1311 => x"83388052",
  1312 => x"7183ffe0",
  1313 => x"800c0288",
  1314 => x"050d0402",
  1315 => x"f8050d73",
  1316 => x"8b118480",
  1317 => x"8080f52d",
  1318 => x"70842a70",
  1319 => x"81065151",
  1320 => x"51518152",
  1321 => x"70833870",
  1322 => x"527183ff",
  1323 => x"e0800c02",
  1324 => x"88050d04",
  1325 => x"02f8050d",
  1326 => x"738b1184",
  1327 => x"808080f5",
  1328 => x"2d70852a",
  1329 => x"70810651",
  1330 => x"51515181",
  1331 => x"52708338",
  1332 => x"70527183",
  1333 => x"ffe0800c",
  1334 => x"0288050d",
  1335 => x"0402fc05",
  1336 => x"0d725180",
  1337 => x"0b84120c",
  1338 => x"80710c02",
  1339 => x"84050d04",
  1340 => x"02f4050d",
  1341 => x"74767008",
  1342 => x"53535370",
  1343 => x"8c388412",
  1344 => x"08730c84",
  1345 => x"8080aa8f",
  1346 => x"04841208",
  1347 => x"84120c84",
  1348 => x"12085170",
  1349 => x"8c387108",
  1350 => x"84140c84",
  1351 => x"8080aaa5",
  1352 => x"04710871",
  1353 => x"0c028c05",
  1354 => x"0d0402f0",
  1355 => x"050d7577",
  1356 => x"84120853",
  1357 => x"545470bf",
  1358 => x"38730852",
  1359 => x"71953872",
  1360 => x"740c7284",
  1361 => x"150c7073",
  1362 => x"0c708414",
  1363 => x"0c848080",
  1364 => x"ab980471",
  1365 => x"08730c71",
  1366 => x"84140c71",
  1367 => x"0851708a",
  1368 => x"3872740c",
  1369 => x"848080aa",
  1370 => x"ee047284",
  1371 => x"120c7272",
  1372 => x"0c848080",
  1373 => x"ab980470",
  1374 => x"730c8411",
  1375 => x"0884140c",
  1376 => x"84110852",
  1377 => x"718b3872",
  1378 => x"84150c84",
  1379 => x"8080ab94",
  1380 => x"0472720c",
  1381 => x"7284120c",
  1382 => x"0290050d",
  1383 => x"0402f405",
  1384 => x"0d88bc15",
  1385 => x"705383ff",
  1386 => x"f2d45253",
  1387 => x"848080a9",
  1388 => x"f02d7252",
  1389 => x"83fff2dc",
  1390 => x"51848080",
  1391 => x"aaaa2d02",
  1392 => x"8c050d04",
  1393 => x"02fdb405",
  1394 => x"0d0282d0",
  1395 => x"050883ff",
  1396 => x"e9ec525a",
  1397 => x"848080d1",
  1398 => x"e72d83ff",
  1399 => x"e080087a",
  1400 => x"52568480",
  1401 => x"8099f72d",
  1402 => x"800b83ff",
  1403 => x"e0800881",
  1404 => x"055a5877",
  1405 => x"792581a0",
  1406 => x"38828454",
  1407 => x"0280c805",
  1408 => x"70547853",
  1409 => x"7a525784",
  1410 => x"80809ba7",
  1411 => x"2d83ffe0",
  1412 => x"8008ff2e",
  1413 => x"09810689",
  1414 => x"38805584",
  1415 => x"8080ada3",
  1416 => x"0402a805",
  1417 => x"70557754",
  1418 => x"765383ff",
  1419 => x"e9ec5255",
  1420 => x"848080d1",
  1421 => x"fa2d83ff",
  1422 => x"e0800880",
  1423 => x"2e903874",
  1424 => x"51848080",
  1425 => x"a98b2d83",
  1426 => x"ffe08008",
  1427 => x"8d3883ff",
  1428 => x"e0800855",
  1429 => x"848080ad",
  1430 => x"a30402bc",
  1431 => x"05848080",
  1432 => x"80e02d70",
  1433 => x"882b83fe",
  1434 => x"80067188",
  1435 => x"2a070288",
  1436 => x"0580c205",
  1437 => x"84808080",
  1438 => x"e02d7088",
  1439 => x"2b83fe80",
  1440 => x"0671882a",
  1441 => x"07728480",
  1442 => x"80290581",
  1443 => x"1c5c5957",
  1444 => x"51578480",
  1445 => x"80abf304",
  1446 => x"0282d405",
  1447 => x"0876710c",
  1448 => x"55815574",
  1449 => x"83ffe080",
  1450 => x"0c0282cc",
  1451 => x"050d0402",
  1452 => x"ffb8050d",
  1453 => x"83fff2dc",
  1454 => x"08705a56",
  1455 => x"75802e83",
  1456 => x"c8387552",
  1457 => x"83fff2dc",
  1458 => x"51848080",
  1459 => x"a9f02d75",
  1460 => x"5283fff2",
  1461 => x"d4518480",
  1462 => x"80aaaa2d",
  1463 => x"f7c41659",
  1464 => x"78802e83",
  1465 => x"a438f7d8",
  1466 => x"165a8284",
  1467 => x"53805279",
  1468 => x"51848080",
  1469 => x"e0f82df9",
  1470 => x"dc165882",
  1471 => x"84538052",
  1472 => x"77518480",
  1473 => x"80e0f82d",
  1474 => x"82845577",
  1475 => x"54828453",
  1476 => x"79526351",
  1477 => x"8480809d",
  1478 => x"b32d83ff",
  1479 => x"e08008ff",
  1480 => x"2e82ee38",
  1481 => x"83fff2d4",
  1482 => x"08577680",
  1483 => x"2ebd38f7",
  1484 => x"c4175675",
  1485 => x"792eaa38",
  1486 => x"7952f7d8",
  1487 => x"17518480",
  1488 => x"80a0ca2d",
  1489 => x"83ffe080",
  1490 => x"08802e95",
  1491 => x"387752f9",
  1492 => x"dc175184",
  1493 => x"8080a0ca",
  1494 => x"2d83ffe0",
  1495 => x"800882b1",
  1496 => x"38841708",
  1497 => x"57848080",
  1498 => x"aeaa0494",
  1499 => x"19848080",
  1500 => x"80f52d56",
  1501 => x"75993883",
  1502 => x"ffe9ec51",
  1503 => x"848080d1",
  1504 => x"e72d83ff",
  1505 => x"e0800879",
  1506 => x"0c848080",
  1507 => x"afb50478",
  1508 => x"52941951",
  1509 => x"848080ab",
  1510 => x"c42d83ff",
  1511 => x"e0800856",
  1512 => x"83ffe080",
  1513 => x"088f3878",
  1514 => x"51848080",
  1515 => x"ab9d2d84",
  1516 => x"8080b19b",
  1517 => x"0402a805",
  1518 => x"70558298",
  1519 => x"1a547908",
  1520 => x"5383ffe9",
  1521 => x"ec525684",
  1522 => x"8080d1fa",
  1523 => x"2d83ffe0",
  1524 => x"8008802e",
  1525 => x"81bb3875",
  1526 => x"51848080",
  1527 => x"a9b42d83",
  1528 => x"ffe08008",
  1529 => x"802e81a9",
  1530 => x"388b5375",
  1531 => x"52849c19",
  1532 => x"51848080",
  1533 => x"de852d61",
  1534 => x"70882b87",
  1535 => x"fc808006",
  1536 => x"7072982b",
  1537 => x"0772882a",
  1538 => x"83fe8006",
  1539 => x"71077398",
  1540 => x"2a078c1d",
  1541 => x"0c515757",
  1542 => x"800b881a",
  1543 => x"0c02bc05",
  1544 => x"84808080",
  1545 => x"e02d7088",
  1546 => x"2b83fe80",
  1547 => x"0671882a",
  1548 => x"07028805",
  1549 => x"80c20584",
  1550 => x"808080e0",
  1551 => x"2d70882b",
  1552 => x"83fe8006",
  1553 => x"71882a07",
  1554 => x"72848080",
  1555 => x"2905841d",
  1556 => x"0c585158",
  1557 => x"ff0b88b0",
  1558 => x"1a0c800b",
  1559 => x"88b41a0c",
  1560 => x"800b901a",
  1561 => x"0cff0b84",
  1562 => x"a81a0cff",
  1563 => x"0b84ac1a",
  1564 => x"0c785283",
  1565 => x"ffe9ec51",
  1566 => x"848080c4",
  1567 => x"a72d83ff",
  1568 => x"e9ec5184",
  1569 => x"808094ad",
  1570 => x"2d785684",
  1571 => x"8080b19b",
  1572 => x"04785184",
  1573 => x"8080ab9d",
  1574 => x"2d805675",
  1575 => x"83ffe080",
  1576 => x"0c0280c8",
  1577 => x"050d0402",
  1578 => x"d0050d7d",
  1579 => x"7f6283ff",
  1580 => x"e9ec0b84",
  1581 => x"808080f5",
  1582 => x"2d705672",
  1583 => x"555a5c56",
  1584 => x"59848080",
  1585 => x"e3b02d83",
  1586 => x"ffe08008",
  1587 => x"83ffe080",
  1588 => x"08782976",
  1589 => x"71317c11",
  1590 => x"585d5758",
  1591 => x"76752785",
  1592 => x"38767b31",
  1593 => x"5a84a819",
  1594 => x"08567776",
  1595 => x"2e098106",
  1596 => x"8c3884ac",
  1597 => x"19085684",
  1598 => x"8080b385",
  1599 => x"0477802e",
  1600 => x"99388116",
  1601 => x"5577752e",
  1602 => x"0981068e",
  1603 => x"387584ac",
  1604 => x"1a085755",
  1605 => x"848080b2",
  1606 => x"a104800b",
  1607 => x"841a0857",
  1608 => x"55747827",
  1609 => x"80d03802",
  1610 => x"b005fc05",
  1611 => x"54745378",
  1612 => x"5283ffe9",
  1613 => x"ec518480",
  1614 => x"80c4af2d",
  1615 => x"83ffe080",
  1616 => x"08a93875",
  1617 => x"5283ffe9",
  1618 => x"ec518480",
  1619 => x"8094fa2d",
  1620 => x"83ffe080",
  1621 => x"085c83ff",
  1622 => x"e0800854",
  1623 => x"74537852",
  1624 => x"83ffe9ec",
  1625 => x"51848080",
  1626 => x"c4b72d7b",
  1627 => x"81165656",
  1628 => x"848080b2",
  1629 => x"a10475ff",
  1630 => x"2e933875",
  1631 => x"84ac1a0c",
  1632 => x"7784a81a",
  1633 => x"0c75ff2e",
  1634 => x"09810689",
  1635 => x"38805584",
  1636 => x"8080b3c7",
  1637 => x"04755283",
  1638 => x"ffe9ec51",
  1639 => x"848080cc",
  1640 => x"d22d7954",
  1641 => x"7f5383ff",
  1642 => x"e080081b",
  1643 => x"5283ffe9",
  1644 => x"ec518480",
  1645 => x"80cda92d",
  1646 => x"795583ff",
  1647 => x"e0800887",
  1648 => x"3883ffe0",
  1649 => x"80085574",
  1650 => x"83ffe080",
  1651 => x"0c02b005",
  1652 => x"0d0402f8",
  1653 => x"050d83ff",
  1654 => x"f2dc5184",
  1655 => x"8080a9dd",
  1656 => x"2d83fff2",
  1657 => x"d4518480",
  1658 => x"80a9dd2d",
  1659 => x"83ffe9e4",
  1660 => x"5283fff2",
  1661 => x"dc518480",
  1662 => x"80aaaa2d",
  1663 => x"810b83ff",
  1664 => x"e1a00c02",
  1665 => x"88050d04",
  1666 => x"02fc050d",
  1667 => x"83ffeaa8",
  1668 => x"73717084",
  1669 => x"05530c74",
  1670 => x"710c5102",
  1671 => x"84050d04",
  1672 => x"02f4050d",
  1673 => x"83ffe1a0",
  1674 => x"08873884",
  1675 => x"8080b3d2",
  1676 => x"2d7483ff",
  1677 => x"eaa00c75",
  1678 => x"83ffeaa4",
  1679 => x"0c83ffe9",
  1680 => x"ec518480",
  1681 => x"80c4bf2d",
  1682 => x"83ffe080",
  1683 => x"085383ff",
  1684 => x"e0800880",
  1685 => x"2e993883",
  1686 => x"ffe08008",
  1687 => x"52848080",
  1688 => x"e8bc5184",
  1689 => x"808082e3",
  1690 => x"2d848080",
  1691 => x"b4fc0481",
  1692 => x"0b83ffe1",
  1693 => x"a40c83ff",
  1694 => x"e0800853",
  1695 => x"7283ffe0",
  1696 => x"800c028c",
  1697 => x"050d0402",
  1698 => x"f8050d83",
  1699 => x"ffe1a008",
  1700 => x"87388480",
  1701 => x"80b3d22d",
  1702 => x"83ffeaa8",
  1703 => x"08527180",
  1704 => x"2e833871",
  1705 => x"2d83ffe9",
  1706 => x"ec518480",
  1707 => x"8094ad2d",
  1708 => x"83ffeaac",
  1709 => x"08527180",
  1710 => x"2e833871",
  1711 => x"2d028805",
  1712 => x"0d0402e8",
  1713 => x"050d7779",
  1714 => x"56568054",
  1715 => x"83ffe1a0",
  1716 => x"08742e09",
  1717 => x"81068738",
  1718 => x"848080b3",
  1719 => x"d22d7352",
  1720 => x"83ffe1a4",
  1721 => x"08802e82",
  1722 => x"ff387581",
  1723 => x"05097077",
  1724 => x"07802576",
  1725 => x"81050970",
  1726 => x"78078025",
  1727 => x"72077752",
  1728 => x"52545153",
  1729 => x"7282e138",
  1730 => x"73538480",
  1731 => x"80b7e504",
  1732 => x"72157084",
  1733 => x"808080f5",
  1734 => x"2d515271",
  1735 => x"80d72e80",
  1736 => x"e8387180",
  1737 => x"d724ad38",
  1738 => x"7180c22e",
  1739 => x"81b03871",
  1740 => x"80c22494",
  1741 => x"3871ab2e",
  1742 => x"80e33871",
  1743 => x"80c12e80",
  1744 => x"d2388480",
  1745 => x"80b7e204",
  1746 => x"7180d22e",
  1747 => x"b2388480",
  1748 => x"80b7e204",
  1749 => x"7180e22e",
  1750 => x"81843871",
  1751 => x"80e2248d",
  1752 => x"387180e1",
  1753 => x"2ead3884",
  1754 => x"8080b7e2",
  1755 => x"047180f2",
  1756 => x"2e8d3871",
  1757 => x"80f72e91",
  1758 => x"38848080",
  1759 => x"b7e20473",
  1760 => x"81075484",
  1761 => x"8080b7e2",
  1762 => x"0473b207",
  1763 => x"54848080",
  1764 => x"b7e20473",
  1765 => x"a6075484",
  1766 => x"8080b7e2",
  1767 => x"04738106",
  1768 => x"5271802e",
  1769 => x"8b387382",
  1770 => x"07548480",
  1771 => x"80b7e204",
  1772 => x"73812a70",
  1773 => x"81065152",
  1774 => x"71802e8b",
  1775 => x"3873b107",
  1776 => x"54848080",
  1777 => x"b7e20473",
  1778 => x"822a7081",
  1779 => x"06515271",
  1780 => x"802e8f38",
  1781 => x"73a70754",
  1782 => x"848080b7",
  1783 => x"e2047388",
  1784 => x"07548113",
  1785 => x"53745184",
  1786 => x"8080d8fa",
  1787 => x"2d83ffe0",
  1788 => x"80087324",
  1789 => x"fe9a3880",
  1790 => x"7481d906",
  1791 => x"555383ff",
  1792 => x"eaa40873",
  1793 => x"2e098106",
  1794 => x"86387381",
  1795 => x"d9065483",
  1796 => x"ffeaa808",
  1797 => x"5271802e",
  1798 => x"8338712d",
  1799 => x"73810652",
  1800 => x"719a3873",
  1801 => x"852a7081",
  1802 => x"06515272",
  1803 => x"a2387180",
  1804 => x"2e983873",
  1805 => x"86065271",
  1806 => x"802e8f38",
  1807 => x"75518480",
  1808 => x"80adaf2d",
  1809 => x"83ffe080",
  1810 => x"08537280",
  1811 => x"2e8b3873",
  1812 => x"88b81484",
  1813 => x"808081b7",
  1814 => x"2d83ffea",
  1815 => x"ac085271",
  1816 => x"802e8338",
  1817 => x"712d7252",
  1818 => x"7183ffe0",
  1819 => x"800c0298",
  1820 => x"050d0480",
  1821 => x"0b83ffe0",
  1822 => x"800c0402",
  1823 => x"f4050d74",
  1824 => x"5283ffe1",
  1825 => x"a0088738",
  1826 => x"848080b3",
  1827 => x"d22d7180",
  1828 => x"2e80da38",
  1829 => x"83ffeaa8",
  1830 => x"08537280",
  1831 => x"2e833872",
  1832 => x"2d901208",
  1833 => x"802e8638",
  1834 => x"800b9013",
  1835 => x"0c800b88",
  1836 => x"130c800b",
  1837 => x"8c130c80",
  1838 => x"0b84130c",
  1839 => x"ff0b88b0",
  1840 => x"130c800b",
  1841 => x"88b4130c",
  1842 => x"800b9013",
  1843 => x"0c715184",
  1844 => x"8080ab9d",
  1845 => x"2d83ffe9",
  1846 => x"ec518480",
  1847 => x"8094ad2d",
  1848 => x"83ffeaac",
  1849 => x"08527180",
  1850 => x"2e833871",
  1851 => x"2d028c05",
  1852 => x"0d0402d0",
  1853 => x"050d7d61",
  1854 => x"6062295a",
  1855 => x"5a5c805b",
  1856 => x"83ffe1a0",
  1857 => x"087b2e09",
  1858 => x"81068738",
  1859 => x"848080b3",
  1860 => x"d22d7b81",
  1861 => x"0509707d",
  1862 => x"0780257a",
  1863 => x"81050970",
  1864 => x"7c078025",
  1865 => x"72075257",
  1866 => x"5156ff5a",
  1867 => x"7581f238",
  1868 => x"88b81984",
  1869 => x"808080f5",
  1870 => x"2d810655",
  1871 => x"74802e81",
  1872 => x"e0387a5a",
  1873 => x"77802e81",
  1874 => x"d8388819",
  1875 => x"088c1a08",
  1876 => x"5856ff5a",
  1877 => x"75772781",
  1878 => x"c8387716",
  1879 => x"55767527",
  1880 => x"85387676",
  1881 => x"31587589",
  1882 => x"2a7683ff",
  1883 => x"065b5580",
  1884 => x"782581ab",
  1885 => x"387980c4",
  1886 => x"38777b31",
  1887 => x"5683ff76",
  1888 => x"25ba3875",
  1889 => x"80258538",
  1890 => x"83ff1656",
  1891 => x"75892c54",
  1892 => x"7a1c5374",
  1893 => x"52785184",
  1894 => x"8080b1a7",
  1895 => x"2d83ffe0",
  1896 => x"8008802e",
  1897 => x"80f93883",
  1898 => x"ffe08008",
  1899 => x"892b83ff",
  1900 => x"e0800816",
  1901 => x"56578480",
  1902 => x"80bc8f04",
  1903 => x"88b01908",
  1904 => x"752ea638",
  1905 => x"815484b0",
  1906 => x"19537452",
  1907 => x"78518480",
  1908 => x"80b1a72d",
  1909 => x"83ffe080",
  1910 => x"08802e80",
  1911 => x"c2387488",
  1912 => x"b01a0c80",
  1913 => x"0b88b41a",
  1914 => x"0c84807a",
  1915 => x"31787c31",
  1916 => x"57577577",
  1917 => x"25833875",
  1918 => x"57765379",
  1919 => x"1984b005",
  1920 => x"527a1c51",
  1921 => x"848080de",
  1922 => x"852d8115",
  1923 => x"55805a76",
  1924 => x"1b881a08",
  1925 => x"18881b0c",
  1926 => x"5b777b24",
  1927 => x"fed7387a",
  1928 => x"5a7983ff",
  1929 => x"e0800c02",
  1930 => x"b0050d04",
  1931 => x"02e8050d",
  1932 => x"80029805",
  1933 => x"84808081",
  1934 => x"b72d7754",
  1935 => x"81538152",
  1936 => x"029805fc",
  1937 => x"05518480",
  1938 => x"80b9f22d",
  1939 => x"83ffe080",
  1940 => x"085583ff",
  1941 => x"e0800881",
  1942 => x"2e098106",
  1943 => x"8b380294",
  1944 => x"05848080",
  1945 => x"80f52d55",
  1946 => x"7483ffe0",
  1947 => x"800c0298",
  1948 => x"050d0402",
  1949 => x"e8050d77",
  1950 => x"797b5853",
  1951 => x"55805372",
  1952 => x"722580d4",
  1953 => x"38ff1254",
  1954 => x"72742580",
  1955 => x"cb387551",
  1956 => x"848080bc",
  1957 => x"ac2d800b",
  1958 => x"83ffe080",
  1959 => x"0824a138",
  1960 => x"74135283",
  1961 => x"ffe08008",
  1962 => x"72848080",
  1963 => x"81b72d81",
  1964 => x"135383ff",
  1965 => x"e080088a",
  1966 => x"2e863873",
  1967 => x"7324cf38",
  1968 => x"80732594",
  1969 => x"38721552",
  1970 => x"80728480",
  1971 => x"8081b72d",
  1972 => x"74528480",
  1973 => x"80bdda04",
  1974 => x"80527183",
  1975 => x"ffe0800c",
  1976 => x"0298050d",
  1977 => x"0402e805",
  1978 => x"0d77797b",
  1979 => x"585454ff",
  1980 => x"5583ffe1",
  1981 => x"a0088738",
  1982 => x"848080b3",
  1983 => x"d22d7452",
  1984 => x"73802e81",
  1985 => x"bc387582",
  1986 => x"32708105",
  1987 => x"09707207",
  1988 => x"80255152",
  1989 => x"5272802e",
  1990 => x"87387452",
  1991 => x"7081a238",
  1992 => x"83ffeaa8",
  1993 => x"08517080",
  1994 => x"2e833870",
  1995 => x"2dff0b88",
  1996 => x"b0150c80",
  1997 => x"0b88b415",
  1998 => x"0c759a38",
  1999 => x"7288150c",
  2000 => x"8c140851",
  2001 => x"70732785",
  2002 => x"38708815",
  2003 => x"0c755584",
  2004 => x"8080bfb2",
  2005 => x"0475812e",
  2006 => x"09810680",
  2007 => x"c5388814",
  2008 => x"08518073",
  2009 => x"249b3872",
  2010 => x"11708816",
  2011 => x"0c8c1508",
  2012 => x"53517171",
  2013 => x"27ba3871",
  2014 => x"88150c84",
  2015 => x"8080bfb0",
  2016 => x"04728105",
  2017 => x"09537073",
  2018 => x"278c3880",
  2019 => x"0b88150c",
  2020 => x"848080bf",
  2021 => x"b0047073",
  2022 => x"3188150c",
  2023 => x"848080bf",
  2024 => x"b0047582",
  2025 => x"2e098106",
  2026 => x"89388c14",
  2027 => x"0888150c",
  2028 => x"805583ff",
  2029 => x"eaac0851",
  2030 => x"70802e83",
  2031 => x"38702d74",
  2032 => x"527183ff",
  2033 => x"e0800c02",
  2034 => x"98050d04",
  2035 => x"02f8050d",
  2036 => x"7352ff51",
  2037 => x"71802ea4",
  2038 => x"3883ffea",
  2039 => x"a8085170",
  2040 => x"802e8338",
  2041 => x"702d7488",
  2042 => x"1308710c",
  2043 => x"5183ffea",
  2044 => x"ac085170",
  2045 => x"802e8338",
  2046 => x"702d8051",
  2047 => x"7083ffe0",
  2048 => x"800c0288",
  2049 => x"050d0402",
  2050 => x"f0050d80",
  2051 => x"54029005",
  2052 => x"fc055275",
  2053 => x"51848080",
  2054 => x"bfcc2d73",
  2055 => x"83ffe080",
  2056 => x"0c029005",
  2057 => x"0d0402f8",
  2058 => x"050d7352",
  2059 => x"ff517180",
  2060 => x"2eb13883",
  2061 => x"ffeaa808",
  2062 => x"5170802e",
  2063 => x"8338702d",
  2064 => x"8812088c",
  2065 => x"13083270",
  2066 => x"81050970",
  2067 => x"72079f2a",
  2068 => x"ff1183ff",
  2069 => x"eaac0854",
  2070 => x"51515252",
  2071 => x"71802e83",
  2072 => x"38712d70",
  2073 => x"83ffe080",
  2074 => x"0c028805",
  2075 => x"0d04800b",
  2076 => x"83ffe080",
  2077 => x"0c0402e4",
  2078 => x"050d787a",
  2079 => x"5755ff57",
  2080 => x"83ffe1a0",
  2081 => x"08873884",
  2082 => x"8080b3d2",
  2083 => x"2d83ffea",
  2084 => x"a8085473",
  2085 => x"802e8338",
  2086 => x"732d7451",
  2087 => x"84808099",
  2088 => x"f72d83ff",
  2089 => x"e08008ff",
  2090 => x"2e098106",
  2091 => x"983883ff",
  2092 => x"e9ec5184",
  2093 => x"8080d1e7",
  2094 => x"2d83ffe0",
  2095 => x"80085784",
  2096 => x"8080c1dc",
  2097 => x"04029c05",
  2098 => x"fc055274",
  2099 => x"51848080",
  2100 => x"abc42d83",
  2101 => x"ffe08008",
  2102 => x"802e9038",
  2103 => x"76537552",
  2104 => x"83ffe9ec",
  2105 => x"51848080",
  2106 => x"d4c92d83",
  2107 => x"ffeaac08",
  2108 => x"5473802e",
  2109 => x"8338732d",
  2110 => x"755476ff",
  2111 => x"2e098106",
  2112 => x"83388054",
  2113 => x"7383ffe0",
  2114 => x"800c029c",
  2115 => x"050d0402",
  2116 => x"ec050d83",
  2117 => x"ffe1a008",
  2118 => x"87388480",
  2119 => x"80b3d22d",
  2120 => x"83ffeaa8",
  2121 => x"08547380",
  2122 => x"2e833873",
  2123 => x"2d775376",
  2124 => x"5283ffe9",
  2125 => x"ec518480",
  2126 => x"80d4e52d",
  2127 => x"83ffe080",
  2128 => x"0883ffea",
  2129 => x"ac085555",
  2130 => x"73802e83",
  2131 => x"38732d74",
  2132 => x"83ffe080",
  2133 => x"0c029405",
  2134 => x"0d0402fd",
  2135 => x"cc050d83",
  2136 => x"ffe1a008",
  2137 => x"87388480",
  2138 => x"80b3d22d",
  2139 => x"83ffeaa8",
  2140 => x"08547380",
  2141 => x"2e833873",
  2142 => x"2d0282a8",
  2143 => x"05705302",
  2144 => x"82bc0508",
  2145 => x"52568480",
  2146 => x"80c0f62d",
  2147 => x"83ffe080",
  2148 => x"08802e80",
  2149 => x"d5388480",
  2150 => x"80c3d404",
  2151 => x"02829c05",
  2152 => x"84808080",
  2153 => x"f52d5473",
  2154 => x"802e9538",
  2155 => x"74528480",
  2156 => x"80e8f051",
  2157 => x"84808082",
  2158 => x"e32d8480",
  2159 => x"80c3d404",
  2160 => x"0282a405",
  2161 => x"08537452",
  2162 => x"848080e8",
  2163 => x"fc518480",
  2164 => x"8082e32d",
  2165 => x"02980570",
  2166 => x"53765255",
  2167 => x"848080c2",
  2168 => x"8f2d83ff",
  2169 => x"e08008ff",
  2170 => x"b33883ff",
  2171 => x"eaac0854",
  2172 => x"73802e83",
  2173 => x"38732d02",
  2174 => x"82b4050d",
  2175 => x"0402e405",
  2176 => x"0d8002a0",
  2177 => x"05f40553",
  2178 => x"79525384",
  2179 => x"8080c0f6",
  2180 => x"2d83ffe0",
  2181 => x"8008732e",
  2182 => x"83388153",
  2183 => x"7283ffe0",
  2184 => x"800c029c",
  2185 => x"050d0481",
  2186 => x"0b83ffe0",
  2187 => x"800c0480",
  2188 => x"0b83ffe0",
  2189 => x"800c0481",
  2190 => x"0b83ffe0",
  2191 => x"800c0402",
  2192 => x"ffb8050d",
  2193 => x"63578058",
  2194 => x"ff0b84c4",
  2195 => x"180c7784",
  2196 => x"c8180c77",
  2197 => x"a4180c76",
  2198 => x"51848080",
  2199 => x"91a52db4",
  2200 => x"170854ff",
  2201 => x"5573782e",
  2202 => x"87dc3881",
  2203 => x"5380c417",
  2204 => x"70537852",
  2205 => x"59732d83",
  2206 => x"ffe08008",
  2207 => x"782e87c6",
  2208 => x"3884c217",
  2209 => x"84808080",
  2210 => x"e02d54fd",
  2211 => x"557381ab",
  2212 => x"aa2e0981",
  2213 => x"0687af38",
  2214 => x"84c31784",
  2215 => x"808080f5",
  2216 => x"2d84c218",
  2217 => x"84808080",
  2218 => x"f52d7182",
  2219 => x"80290555",
  2220 => x"55fc5573",
  2221 => x"82d4d52e",
  2222 => x"09810687",
  2223 => x"89388486",
  2224 => x"17848080",
  2225 => x"80f52d70",
  2226 => x"81ff0655",
  2227 => x"56738f26",
  2228 => x"a0388174",
  2229 => x"2b7083b0",
  2230 => x"e0065555",
  2231 => x"73782e09",
  2232 => x"81069938",
  2233 => x"74810654",
  2234 => x"73782e09",
  2235 => x"810680d0",
  2236 => x"387581ff",
  2237 => x"06547386",
  2238 => x"2680c538",
  2239 => x"848d1784",
  2240 => x"808080f5",
  2241 => x"2d848c18",
  2242 => x"84808080",
  2243 => x"f52d7181",
  2244 => x"800a2971",
  2245 => x"84808029",
  2246 => x"05848b1a",
  2247 => x"84808080",
  2248 => x"f52d7082",
  2249 => x"80291284",
  2250 => x"8a1c8480",
  2251 => x"8080f52d",
  2252 => x"5574059c",
  2253 => x"1c0c5956",
  2254 => x"56588480",
  2255 => x"80c6c404",
  2256 => x"779c180c",
  2257 => x"81537852",
  2258 => x"9c170851",
  2259 => x"b4170854",
  2260 => x"732dff55",
  2261 => x"83ffe080",
  2262 => x"08802e85",
  2263 => x"e93880d0",
  2264 => x"17848080",
  2265 => x"80f52d80",
  2266 => x"cf188480",
  2267 => x"8080f52d",
  2268 => x"7072882b",
  2269 => x"0756415f",
  2270 => x"fe557384",
  2271 => x"802e0981",
  2272 => x"0685c338",
  2273 => x"80d11784",
  2274 => x"808080f5",
  2275 => x"2d778480",
  2276 => x"8081b72d",
  2277 => x"80d31784",
  2278 => x"808080f5",
  2279 => x"2d80d218",
  2280 => x"84808080",
  2281 => x"f52d7072",
  2282 => x"882b0780",
  2283 => x"d41a8480",
  2284 => x"8080f52d",
  2285 => x"7081ff06",
  2286 => x"80d61c84",
  2287 => x"808080f5",
  2288 => x"2d80d51d",
  2289 => x"84808080",
  2290 => x"f52d7072",
  2291 => x"882b075b",
  2292 => x"415f5a41",
  2293 => x"5b434173",
  2294 => x"a8188480",
  2295 => x"80818a2d",
  2296 => x"80db1784",
  2297 => x"808080f5",
  2298 => x"2d80da18",
  2299 => x"84808080",
  2300 => x"f52d7072",
  2301 => x"882b0756",
  2302 => x"5e5c7380",
  2303 => x"2e8b3873",
  2304 => x"a0180c84",
  2305 => x"8080c8c7",
  2306 => x"0480eb17",
  2307 => x"84808080",
  2308 => x"f52d80ea",
  2309 => x"18848080",
  2310 => x"80f52d71",
  2311 => x"81800a29",
  2312 => x"71848080",
  2313 => x"290580e9",
  2314 => x"1a848080",
  2315 => x"80f52d70",
  2316 => x"82802912",
  2317 => x"80e81c84",
  2318 => x"808080f5",
  2319 => x"2d547305",
  2320 => x"a01c0c53",
  2321 => x"56595580",
  2322 => x"f3178480",
  2323 => x"8080f52d",
  2324 => x"80f21884",
  2325 => x"808080f5",
  2326 => x"2d718180",
  2327 => x"0a297184",
  2328 => x"80802905",
  2329 => x"80f11a84",
  2330 => x"808080f5",
  2331 => x"2d708280",
  2332 => x"291280f0",
  2333 => x"1c848080",
  2334 => x"80f52d54",
  2335 => x"7305881c",
  2336 => x"0c80f51b",
  2337 => x"84808080",
  2338 => x"f52d80f4",
  2339 => x"1c848080",
  2340 => x"80f52d71",
  2341 => x"82802905",
  2342 => x"53515356",
  2343 => x"59557398",
  2344 => x"18848080",
  2345 => x"818a2d75",
  2346 => x"a0180829",
  2347 => x"701a8c19",
  2348 => x"0ca81884",
  2349 => x"808080e0",
  2350 => x"2d70852b",
  2351 => x"83ff1152",
  2352 => x"58555873",
  2353 => x"80258538",
  2354 => x"87fe1654",
  2355 => x"73892a90",
  2356 => x"180c9c17",
  2357 => x"08197094",
  2358 => x"190c7805",
  2359 => x"84180c84",
  2360 => x"c3178480",
  2361 => x"8080f52d",
  2362 => x"84c21884",
  2363 => x"808080f5",
  2364 => x"2d718280",
  2365 => x"29055555",
  2366 => x"fd557382",
  2367 => x"d4d52e09",
  2368 => x"810682c2",
  2369 => x"3879882b",
  2370 => x"83fe8006",
  2371 => x"7b81ff06",
  2372 => x"7012852b",
  2373 => x"61882b83",
  2374 => x"fe800663",
  2375 => x"81ff0671",
  2376 => x"05705751",
  2377 => x"527105ff",
  2378 => x"05535556",
  2379 => x"848080e2",
  2380 => x"dd2d83ff",
  2381 => x"e080087c",
  2382 => x"882b83fe",
  2383 => x"80067e81",
  2384 => x"ff067105",
  2385 => x"705c5155",
  2386 => x"5a73bd38",
  2387 => x"80eb1784",
  2388 => x"808080f5",
  2389 => x"2d80ea18",
  2390 => x"84808080",
  2391 => x"f52d7181",
  2392 => x"800a2971",
  2393 => x"84808029",
  2394 => x"0580e91a",
  2395 => x"84808080",
  2396 => x"f52d7082",
  2397 => x"80291280",
  2398 => x"e81c8480",
  2399 => x"8080f52d",
  2400 => x"5574055d",
  2401 => x"59565658",
  2402 => x"80d81784",
  2403 => x"808080f5",
  2404 => x"2d80d718",
  2405 => x"84808080",
  2406 => x"f52d7182",
  2407 => x"80290570",
  2408 => x"5a555573",
  2409 => x"bd3880e7",
  2410 => x"17848080",
  2411 => x"80f52d80",
  2412 => x"e6188480",
  2413 => x"8080f52d",
  2414 => x"7181800a",
  2415 => x"29718480",
  2416 => x"80290580",
  2417 => x"e51a8480",
  2418 => x"8080f52d",
  2419 => x"70828029",
  2420 => x"1280e41c",
  2421 => x"84808080",
  2422 => x"f52d5473",
  2423 => x"05545956",
  2424 => x"56586088",
  2425 => x"2b83fe80",
  2426 => x"066281ff",
  2427 => x"067f81ff",
  2428 => x"06577105",
  2429 => x"767b2905",
  2430 => x"7971317c",
  2431 => x"31798480",
  2432 => x"8080f52d",
  2433 => x"52585154",
  2434 => x"fb557380",
  2435 => x"2eb83873",
  2436 => x"52755184",
  2437 => x"8080e3b0",
  2438 => x"2d9ff40b",
  2439 => x"83ffe080",
  2440 => x"0827a338",
  2441 => x"83ffe080",
  2442 => x"0883fff4",
  2443 => x"26913880",
  2444 => x"0b88180c",
  2445 => x"800bb018",
  2446 => x"0c848080",
  2447 => x"ccc40481",
  2448 => x"0bb0180c",
  2449 => x"80557483",
  2450 => x"ffe0800c",
  2451 => x"0280c805",
  2452 => x"0d0402e8",
  2453 => x"050d7779",
  2454 => x"5755b015",
  2455 => x"08af38a8",
  2456 => x"15848080",
  2457 => x"80e02d53",
  2458 => x"72802584",
  2459 => x"388f1353",
  2460 => x"72842a84",
  2461 => x"16080575",
  2462 => x"84808080",
  2463 => x"f52dfe18",
  2464 => x"71297205",
  2465 => x"52565484",
  2466 => x"8080cd9e",
  2467 => x"04748480",
  2468 => x"8080f52d",
  2469 => x"fe177129",
  2470 => x"84170805",
  2471 => x"51547383",
  2472 => x"ffe0800c",
  2473 => x"0298050d",
  2474 => x"0402f005",
  2475 => x"0d785377",
  2476 => x"52765175",
  2477 => x"b4110851",
  2478 => x"54732d02",
  2479 => x"90050d04",
  2480 => x"02f0050d",
  2481 => x"78537752",
  2482 => x"765175b8",
  2483 => x"11085154",
  2484 => x"732d0290",
  2485 => x"050d0402",
  2486 => x"d4050d7c",
  2487 => x"7e60625e",
  2488 => x"5c565780",
  2489 => x"705559b0",
  2490 => x"1708792e",
  2491 => x"09810683",
  2492 => x"38815478",
  2493 => x"5874a138",
  2494 => x"73587380",
  2495 => x"2e9a3878",
  2496 => x"55799018",
  2497 => x"082781a0",
  2498 => x"389c1708",
  2499 => x"8c180805",
  2500 => x"1a548480",
  2501 => x"80cef604",
  2502 => x"74778480",
  2503 => x"8080f52d",
  2504 => x"70547b53",
  2505 => x"55568480",
  2506 => x"80e3b02d",
  2507 => x"83ffe080",
  2508 => x"0874297a",
  2509 => x"71315a54",
  2510 => x"7783ffe0",
  2511 => x"8008279d",
  2512 => x"3883ffe0",
  2513 => x"80085475",
  2514 => x"52765184",
  2515 => x"808094fa",
  2516 => x"2d83ffe0",
  2517 => x"8008ff15",
  2518 => x"555673eb",
  2519 => x"38805575",
  2520 => x"ff2e80c4",
  2521 => x"38755276",
  2522 => x"51848080",
  2523 => x"ccd22d83",
  2524 => x"ffe08008",
  2525 => x"19547a80",
  2526 => x"2e8b3881",
  2527 => x"537a5284",
  2528 => x"8080cf9a",
  2529 => x"04815573",
  2530 => x"84c41808",
  2531 => x"2e9a3873",
  2532 => x"84c4180c",
  2533 => x"745380c4",
  2534 => x"17527351",
  2535 => x"b4170854",
  2536 => x"732d83ff",
  2537 => x"e0800855",
  2538 => x"7483ffe0",
  2539 => x"800c02ac",
  2540 => x"050d0402",
  2541 => x"d8050d7b",
  2542 => x"7d7f61b0",
  2543 => x"14087081",
  2544 => x"0509b016",
  2545 => x"08710770",
  2546 => x"09709f2a",
  2547 => x"51515151",
  2548 => x"585c5c59",
  2549 => x"5677bf38",
  2550 => x"81707506",
  2551 => x"55577380",
  2552 => x"2eb43877",
  2553 => x"54799017",
  2554 => x"082780f4",
  2555 => x"389c1608",
  2556 => x"8c170805",
  2557 => x"1ab41708",
  2558 => x"56547880",
  2559 => x"2e8b3876",
  2560 => x"53785284",
  2561 => x"8080d0d6",
  2562 => x"047384c4",
  2563 => x"170c7653",
  2564 => x"848080d0",
  2565 => x"d204b416",
  2566 => x"08557880",
  2567 => x"2e9c3877",
  2568 => x"52755184",
  2569 => x"8080ccd2",
  2570 => x"2d815378",
  2571 => x"5283ffe0",
  2572 => x"80081a51",
  2573 => x"848080d0",
  2574 => x"d8047752",
  2575 => x"75518480",
  2576 => x"80ccd22d",
  2577 => x"83ffe080",
  2578 => x"081a7084",
  2579 => x"c4180c54",
  2580 => x"815380c4",
  2581 => x"16527351",
  2582 => x"742d83ff",
  2583 => x"e0800854",
  2584 => x"7383ffe0",
  2585 => x"800c02a8",
  2586 => x"050d0402",
  2587 => x"f0050d75",
  2588 => x"848080e9",
  2589 => x"8c525484",
  2590 => x"808082e3",
  2591 => x"2d848080",
  2592 => x"e99c53b0",
  2593 => x"1408812e",
  2594 => x"87388480",
  2595 => x"80e9a453",
  2596 => x"72528480",
  2597 => x"80e9ac51",
  2598 => x"84808082",
  2599 => x"e32d8814",
  2600 => x"08528480",
  2601 => x"80e9b851",
  2602 => x"84808082",
  2603 => x"e32d9414",
  2604 => x"08528480",
  2605 => x"80e9d851",
  2606 => x"84808082",
  2607 => x"e32d8414",
  2608 => x"08528480",
  2609 => x"80e9f051",
  2610 => x"84808082",
  2611 => x"e32d7384",
  2612 => x"808080f5",
  2613 => x"2d528480",
  2614 => x"80ea8c51",
  2615 => x"84808082",
  2616 => x"e32d0290",
  2617 => x"050d0402",
  2618 => x"fc050d72",
  2619 => x"88110883",
  2620 => x"ffe0800c",
  2621 => x"51028405",
  2622 => x"0d0402ff",
  2623 => x"ac050d66",
  2624 => x"686a4141",
  2625 => x"5e805d81",
  2626 => x"520280d4",
  2627 => x"05ec0551",
  2628 => x"848080a8",
  2629 => x"8b2d8054",
  2630 => x"7c53811d",
  2631 => x"60537e52",
  2632 => x"5d848080",
  2633 => x"cdd72d83",
  2634 => x"ffe08008",
  2635 => x"802e828b",
  2636 => x"38805b7a",
  2637 => x"a0291e80",
  2638 => x"c4057052",
  2639 => x"58848080",
  2640 => x"a8c72d83",
  2641 => x"ffe08008",
  2642 => x"802e81db",
  2643 => x"380280c4",
  2644 => x"05598d53",
  2645 => x"80527851",
  2646 => x"848080e0",
  2647 => x"f82d8057",
  2648 => x"76197719",
  2649 => x"57557584",
  2650 => x"808080f5",
  2651 => x"2d758480",
  2652 => x"8081b72d",
  2653 => x"81177081",
  2654 => x"ff065855",
  2655 => x"877727e0",
  2656 => x"38805a88",
  2657 => x"02840580",
  2658 => x"c5055d57",
  2659 => x"761c7719",
  2660 => x"56567484",
  2661 => x"808080f5",
  2662 => x"2d768480",
  2663 => x"8081b72d",
  2664 => x"74848080",
  2665 => x"80f52d55",
  2666 => x"74a02e83",
  2667 => x"38815a81",
  2668 => x"177081ff",
  2669 => x"0658558a",
  2670 => x"7727d138",
  2671 => x"79802ea2",
  2672 => x"380280c4",
  2673 => x"05848080",
  2674 => x"80f52d55",
  2675 => x"74ae2e92",
  2676 => x"38ae0280",
  2677 => x"d0058480",
  2678 => x"8081b72d",
  2679 => x"848080d3",
  2680 => x"ed04a002",
  2681 => x"80d00584",
  2682 => x"808081b7",
  2683 => x"2d7e5278",
  2684 => x"51848080",
  2685 => x"a0ca2d83",
  2686 => x"ffe08008",
  2687 => x"802e9538",
  2688 => x"a0537752",
  2689 => x"69518480",
  2690 => x"80de852d",
  2691 => x"81558480",
  2692 => x"80d4bd04",
  2693 => x"83ffe080",
  2694 => x"08520280",
  2695 => x"d405ec05",
  2696 => x"51848080",
  2697 => x"a88b2d81",
  2698 => x"1b7081ff",
  2699 => x"065c558f",
  2700 => x"7b27fdff",
  2701 => x"38848080",
  2702 => x"d2960480",
  2703 => x"557483ff",
  2704 => x"e0800c02",
  2705 => x"80d4050d",
  2706 => x"0402fc05",
  2707 => x"0d737584",
  2708 => x"120c5180",
  2709 => x"710c800b",
  2710 => x"88128480",
  2711 => x"8081b72d",
  2712 => x"0284050d",
  2713 => x"0402ffb4",
  2714 => x"050d6466",
  2715 => x"68405b56",
  2716 => x"80520280",
  2717 => x"cc05ec05",
  2718 => x"51848080",
  2719 => x"a88b2d80",
  2720 => x"54790853",
  2721 => x"841a0852",
  2722 => x"75518480",
  2723 => x"80cdd72d",
  2724 => x"83ffe080",
  2725 => x"08802e83",
  2726 => x"d338881a",
  2727 => x"84808080",
  2728 => x"f52d5978",
  2729 => x"8f2683ae",
  2730 => x"3878a029",
  2731 => x"1680c405",
  2732 => x"70525884",
  2733 => x"8080a8c7",
  2734 => x"2d83ffe0",
  2735 => x"8008802e",
  2736 => x"83863880",
  2737 => x"520280cc",
  2738 => x"05ec0551",
  2739 => x"848080a8",
  2740 => x"8b2d02bc",
  2741 => x"055b8d53",
  2742 => x"80527a51",
  2743 => x"848080e0",
  2744 => x"f82d8057",
  2745 => x"761b7719",
  2746 => x"57557584",
  2747 => x"808080f5",
  2748 => x"2d758480",
  2749 => x"8081b72d",
  2750 => x"81177081",
  2751 => x"ff065855",
  2752 => x"877727e0",
  2753 => x"38805c88",
  2754 => x"028405bd",
  2755 => x"055e5776",
  2756 => x"1d771956",
  2757 => x"56748480",
  2758 => x"8080f52d",
  2759 => x"76848080",
  2760 => x"81b72d74",
  2761 => x"84808080",
  2762 => x"f52d5574",
  2763 => x"a02e8338",
  2764 => x"815c8117",
  2765 => x"7081ff06",
  2766 => x"58558a77",
  2767 => x"27d1387b",
  2768 => x"802ea138",
  2769 => x"02bc0584",
  2770 => x"808080f5",
  2771 => x"2d5574ae",
  2772 => x"2e9238ae",
  2773 => x"0280c805",
  2774 => x"84808081",
  2775 => x"b72d8480",
  2776 => x"80d6ef04",
  2777 => x"a00280c8",
  2778 => x"05848080",
  2779 => x"81b72d7a",
  2780 => x"527d5184",
  2781 => x"8080a482",
  2782 => x"2d775184",
  2783 => x"8080a98b",
  2784 => x"2d83ffe0",
  2785 => x"8008802e",
  2786 => x"9238810b",
  2787 => x"82841f84",
  2788 => x"808081b7",
  2789 => x"2d848080",
  2790 => x"d7a90483",
  2791 => x"ffe08008",
  2792 => x"82841f84",
  2793 => x"808081b7",
  2794 => x"2d9c1884",
  2795 => x"808080f5",
  2796 => x"2d9d1984",
  2797 => x"808080f5",
  2798 => x"2d71982b",
  2799 => x"71902b07",
  2800 => x"9e1b8480",
  2801 => x"8080f52d",
  2802 => x"70882b72",
  2803 => x"079f1d84",
  2804 => x"808080f5",
  2805 => x"2d710770",
  2806 => x"882b87fc",
  2807 => x"80800670",
  2808 => x"72982b07",
  2809 => x"72882a83",
  2810 => x"fe800671",
  2811 => x"0773982a",
  2812 => x"0766828c",
  2813 => x"050c5153",
  2814 => x"51525957",
  2815 => x"951a8480",
  2816 => x"8080f52d",
  2817 => x"941b8480",
  2818 => x"8080f52d",
  2819 => x"71982b71",
  2820 => x"902b079b",
  2821 => x"1d848080",
  2822 => x"80f52d9a",
  2823 => x"1e848080",
  2824 => x"80f52d71",
  2825 => x"882b0772",
  2826 => x"07648288",
  2827 => x"050c811f",
  2828 => x"53555a58",
  2829 => x"515c5774",
  2830 => x"881b8480",
  2831 => x"8081b72d",
  2832 => x"81558480",
  2833 => x"80d8ee04",
  2834 => x"81197081",
  2835 => x"ff065a55",
  2836 => x"848080d5",
  2837 => x"a3047908",
  2838 => x"81057a0c",
  2839 => x"800b881b",
  2840 => x"84808081",
  2841 => x"b72d8480",
  2842 => x"80d4ff04",
  2843 => x"80557483",
  2844 => x"ffe0800c",
  2845 => x"0280cc05",
  2846 => x"0d0402f4",
  2847 => x"050d7452",
  2848 => x"80727081",
  2849 => x"05548480",
  2850 => x"8080f52d",
  2851 => x"52537073",
  2852 => x"2e933881",
  2853 => x"13727081",
  2854 => x"05548480",
  2855 => x"8080f52d",
  2856 => x"525370ef",
  2857 => x"387283ff",
  2858 => x"e0800c02",
  2859 => x"8c050d04",
  2860 => x"02f0050d",
  2861 => x"75777156",
  2862 => x"54527270",
  2863 => x"81055484",
  2864 => x"808080f5",
  2865 => x"2d517072",
  2866 => x"70810554",
  2867 => x"84808081",
  2868 => x"b72d70e6",
  2869 => x"387383ff",
  2870 => x"e0800c02",
  2871 => x"90050d04",
  2872 => x"02e4050d",
  2873 => x"787a7c72",
  2874 => x"5a545553",
  2875 => x"848080da",
  2876 => x"81048114",
  2877 => x"54747370",
  2878 => x"81055584",
  2879 => x"808081b7",
  2880 => x"2d807484",
  2881 => x"808080f5",
  2882 => x"2d7081ff",
  2883 => x"06535656",
  2884 => x"70762e83",
  2885 => x"38815671",
  2886 => x"81050970",
  2887 => x"73079f2a",
  2888 => x"707806ff",
  2889 => x"15555151",
  2890 => x"5170c738",
  2891 => x"71ff2e96",
  2892 => x"38807370",
  2893 => x"81055584",
  2894 => x"808081b7",
  2895 => x"2dff1252",
  2896 => x"848080da",
  2897 => x"ac047683",
  2898 => x"ffe0800c",
  2899 => x"029c050d",
  2900 => x"0402f005",
  2901 => x"0d757771",
  2902 => x"56545271",
  2903 => x"70810553",
  2904 => x"84808080",
  2905 => x"f52d5170",
  2906 => x"f2387270",
  2907 => x"81055484",
  2908 => x"808080f5",
  2909 => x"2d517072",
  2910 => x"70810554",
  2911 => x"84808081",
  2912 => x"b72d70e6",
  2913 => x"387383ff",
  2914 => x"e0800c02",
  2915 => x"90050d04",
  2916 => x"02ec050d",
  2917 => x"76787a72",
  2918 => x"58555552",
  2919 => x"71708105",
  2920 => x"53848080",
  2921 => x"80f52d51",
  2922 => x"70f23884",
  2923 => x"8080dbbf",
  2924 => x"04ff1353",
  2925 => x"72ff2e9a",
  2926 => x"38811281",
  2927 => x"15555273",
  2928 => x"84808080",
  2929 => x"f52d5170",
  2930 => x"72848080",
  2931 => x"81b72d70",
  2932 => x"e0388072",
  2933 => x"84808081",
  2934 => x"b72d7483",
  2935 => x"ffe0800c",
  2936 => x"0294050d",
  2937 => x"0402f005",
  2938 => x"0d757752",
  2939 => x"52848080",
  2940 => x"dc890470",
  2941 => x"84808080",
  2942 => x"f52d5472",
  2943 => x"742e0981",
  2944 => x"06923881",
  2945 => x"12811252",
  2946 => x"52718480",
  2947 => x"8080f52d",
  2948 => x"5372e038",
  2949 => x"71848080",
  2950 => x"80f52d71",
  2951 => x"84808080",
  2952 => x"f52d7171",
  2953 => x"3183ffe0",
  2954 => x"800c5252",
  2955 => x"0290050d",
  2956 => x"0402ec05",
  2957 => x"0d76787a",
  2958 => x"70555354",
  2959 => x"5470802e",
  2960 => x"80c33884",
  2961 => x"8080dcd7",
  2962 => x"04ff1151",
  2963 => x"70802ea1",
  2964 => x"38811481",
  2965 => x"14545473",
  2966 => x"84808080",
  2967 => x"f52d5271",
  2968 => x"802e8e38",
  2969 => x"72848080",
  2970 => x"80f52d55",
  2971 => x"71752ed9",
  2972 => x"38738480",
  2973 => x"8080f52d",
  2974 => x"73848080",
  2975 => x"80f52d71",
  2976 => x"71315454",
  2977 => x"547183ff",
  2978 => x"e0800c02",
  2979 => x"94050d04",
  2980 => x"02f4050d",
  2981 => x"74765451",
  2982 => x"848080dd",
  2983 => x"a6047173",
  2984 => x"2e8f3881",
  2985 => x"11517084",
  2986 => x"808080f5",
  2987 => x"2d5271ee",
  2988 => x"387083ff",
  2989 => x"e0800c02",
  2990 => x"8c050d04",
  2991 => x"02ec050d",
  2992 => x"76785653",
  2993 => x"80738480",
  2994 => x"8080f52d",
  2995 => x"7081ff06",
  2996 => x"53535470",
  2997 => x"742ea338",
  2998 => x"7181ff06",
  2999 => x"5170752e",
  3000 => x"09810683",
  3001 => x"38725481",
  3002 => x"13708480",
  3003 => x"8080f52d",
  3004 => x"7081ff06",
  3005 => x"53535370",
  3006 => x"df387383",
  3007 => x"ffe0800c",
  3008 => x"0294050d",
  3009 => x"0402e805",
  3010 => x"0d77797b",
  3011 => x"72720783",
  3012 => x"06545456",
  3013 => x"5670802e",
  3014 => x"aa387476",
  3015 => x"5253ff12",
  3016 => x"5271ff2e",
  3017 => x"80f43872",
  3018 => x"70810554",
  3019 => x"84808080",
  3020 => x"f52d7170",
  3021 => x"81055384",
  3022 => x"808081b7",
  3023 => x"2d848080",
  3024 => x"de9e0474",
  3025 => x"7673822a",
  3026 => x"ff055354",
  3027 => x"5470ff2e",
  3028 => x"96387370",
  3029 => x"84055508",
  3030 => x"73708405",
  3031 => x"550cff11",
  3032 => x"51848080",
  3033 => x"decd0471",
  3034 => x"fc067016",
  3035 => x"55760572",
  3036 => x"8306ff05",
  3037 => x"525370ff",
  3038 => x"2ea03873",
  3039 => x"70810555",
  3040 => x"84808080",
  3041 => x"f52d7370",
  3042 => x"81055584",
  3043 => x"808081b7",
  3044 => x"2dff1151",
  3045 => x"848080de",
  3046 => x"f6047583",
  3047 => x"ffe0800c",
  3048 => x"0298050d",
  3049 => x"0402f005",
  3050 => x"0d757078",
  3051 => x"ff1b5454",
  3052 => x"545470ff",
  3053 => x"2ea03871",
  3054 => x"70810553",
  3055 => x"84808080",
  3056 => x"f52d7370",
  3057 => x"81055584",
  3058 => x"808081b7",
  3059 => x"2dff1151",
  3060 => x"848080df",
  3061 => x"b2047383",
  3062 => x"ffe0800c",
  3063 => x"0290050d",
  3064 => x"0402ec05",
  3065 => x"0d787779",
  3066 => x"53545284",
  3067 => x"8080dfff",
  3068 => x"04ff1252",
  3069 => x"71ff2e9c",
  3070 => x"38811381",
  3071 => x"12525370",
  3072 => x"84808080",
  3073 => x"f52d7384",
  3074 => x"808080f5",
  3075 => x"2d565473",
  3076 => x"752ede38",
  3077 => x"72848080",
  3078 => x"80f52d71",
  3079 => x"84808080",
  3080 => x"f52d7171",
  3081 => x"3183ffe0",
  3082 => x"800c5253",
  3083 => x"0294050d",
  3084 => x"0402f005",
  3085 => x"0d767877",
  3086 => x"54525384",
  3087 => x"8080e0cc",
  3088 => x"04ff1151",
  3089 => x"70ff2e94",
  3090 => x"38811252",
  3091 => x"71848080",
  3092 => x"80f52d54",
  3093 => x"72742e09",
  3094 => x"8106e638",
  3095 => x"71728480",
  3096 => x"8080f52d",
  3097 => x"53517272",
  3098 => x"2e833880",
  3099 => x"517083ff",
  3100 => x"e0800c02",
  3101 => x"90050d04",
  3102 => x"02f0050d",
  3103 => x"757771ff",
  3104 => x"1b545455",
  3105 => x"5370ff2e",
  3106 => x"96387372",
  3107 => x"70810554",
  3108 => x"84808081",
  3109 => x"b72dff11",
  3110 => x"51848080",
  3111 => x"e1850472",
  3112 => x"83ffe080",
  3113 => x"0c029005",
  3114 => x"0d0402f0",
  3115 => x"050d7552",
  3116 => x"848080e1",
  3117 => x"b9048112",
  3118 => x"52807284",
  3119 => x"808080f5",
  3120 => x"2d7081ff",
  3121 => x"06535454",
  3122 => x"70742e83",
  3123 => x"38815470",
  3124 => x"a02e8438",
  3125 => x"73e03872",
  3126 => x"81ff0651",
  3127 => x"70a02e09",
  3128 => x"81069238",
  3129 => x"81127084",
  3130 => x"808080f5",
  3131 => x"2d525284",
  3132 => x"8080e1dc",
  3133 => x"04718480",
  3134 => x"8080f52d",
  3135 => x"70545170",
  3136 => x"802e8338",
  3137 => x"71537283",
  3138 => x"ffe0800c",
  3139 => x"0290050d",
  3140 => x"0402e805",
  3141 => x"0d777957",
  3142 => x"55805473",
  3143 => x"7524b338",
  3144 => x"75742953",
  3145 => x"72752e09",
  3146 => x"81068938",
  3147 => x"80538480",
  3148 => x"80e2d204",
  3149 => x"74732591",
  3150 => x"38737629",
  3151 => x"76317571",
  3152 => x"31515384",
  3153 => x"8080e2d2",
  3154 => x"04811454",
  3155 => x"848080e2",
  3156 => x"9b047283",
  3157 => x"ffe0800c",
  3158 => x"0298050d",
  3159 => x"0402e005",
  3160 => x"0d797b58",
  3161 => x"56807059",
  3162 => x"54775377",
  3163 => x"762eb638",
  3164 => x"77762499",
  3165 => x"38811477",
  3166 => x"19595475",
  3167 => x"7427ea38",
  3168 => x"72547485",
  3169 => x"249f3884",
  3170 => x"8080e3a3",
  3171 => x"04737729",
  3172 => x"77317671",
  3173 => x"31902b70",
  3174 => x"902c5156",
  3175 => x"53848080",
  3176 => x"e3800472",
  3177 => x"547383ff",
  3178 => x"e0800c02",
  3179 => x"a0050d04",
  3180 => x"02f8050d",
  3181 => x"74527351",
  3182 => x"848080e2",
  3183 => x"dd2d0288",
  3184 => x"050d0402",
  3185 => x"f8050d74",
  3186 => x"52735184",
  3187 => x"8080e291",
  3188 => x"2d028805",
  3189 => x"0d0402c0",
  3190 => x"050d8480",
  3191 => x"80eaa851",
  3192 => x"84808082",
  3193 => x"e32d8480",
  3194 => x"80eac051",
  3195 => x"84808082",
  3196 => x"e32d8480",
  3197 => x"80ead851",
  3198 => x"84808082",
  3199 => x"e32d8480",
  3200 => x"8091942d",
  3201 => x"83ffe080",
  3202 => x"08810655",
  3203 => x"7481e838",
  3204 => x"848080ea",
  3205 => x"ec518480",
  3206 => x"8082e32d",
  3207 => x"8480808d",
  3208 => x"bf2d8480",
  3209 => x"80b3d22d",
  3210 => x"84808090",
  3211 => x"e4528480",
  3212 => x"8090b251",
  3213 => x"848080b4",
  3214 => x"a02d83ff",
  3215 => x"e0800880",
  3216 => x"2e80d238",
  3217 => x"848080eb",
  3218 => x"84518480",
  3219 => x"8082e32d",
  3220 => x"81558480",
  3221 => x"80e7b904",
  3222 => x"83ffe080",
  3223 => x"08549080",
  3224 => x"80538152",
  3225 => x"80c0c084",
  3226 => x"51848080",
  3227 => x"b9f22d83",
  3228 => x"ffe08008",
  3229 => x"52848080",
  3230 => x"eba05184",
  3231 => x"808082e3",
  3232 => x"2d745184",
  3233 => x"8080b8fb",
  3234 => x"2d848080",
  3235 => x"b5872d84",
  3236 => x"8080e6aa",
  3237 => x"04848080",
  3238 => x"ebb45184",
  3239 => x"808082e3",
  3240 => x"2d848080",
  3241 => x"ebd05184",
  3242 => x"8080c2da",
  3243 => x"2d848080",
  3244 => x"ebd45184",
  3245 => x"808082e3",
  3246 => x"2d80538e",
  3247 => x"5202b005",
  3248 => x"70525584",
  3249 => x"808086ae",
  3250 => x"2d848080",
  3251 => x"ebe45274",
  3252 => x"51848080",
  3253 => x"b5c22d83",
  3254 => x"ffe08008",
  3255 => x"5583ffe0",
  3256 => x"8008fef4",
  3257 => x"38848080",
  3258 => x"ebe85184",
  3259 => x"808082e3",
  3260 => x"2d848080",
  3261 => x"e5ad0484",
  3262 => x"8080ec84",
  3263 => x"51848080",
  3264 => x"82e32d84",
  3265 => x"808087c6",
  3266 => x"2d805383",
  3267 => x"ffe08008",
  3268 => x"520280c0",
  3269 => x"05e40551",
  3270 => x"84808086",
  3271 => x"ae2d8480",
  3272 => x"80ecb051",
  3273 => x"84808082",
  3274 => x"e32d8059",
  3275 => x"78822b80",
  3276 => x"c0c08711",
  3277 => x"84808080",
  3278 => x"f52d80c0",
  3279 => x"c0861284",
  3280 => x"808080f5",
  3281 => x"2d71982b",
  3282 => x"71902b07",
  3283 => x"80c0c085",
  3284 => x"14848080",
  3285 => x"80f52d70",
  3286 => x"882b7207",
  3287 => x"80c0c084",
  3288 => x"16848080",
  3289 => x"80f52d71",
  3290 => x"0770882a",
  3291 => x"83fe8006",
  3292 => x"7072982a",
  3293 => x"0772882b",
  3294 => x"87fc8080",
  3295 => x"06710773",
  3296 => x"982b0779",
  3297 => x"0c515351",
  3298 => x"52535859",
  3299 => x"57588119",
  3300 => x"5983ffff",
  3301 => x"7925ff94",
  3302 => x"38848080",
  3303 => x"ecb45184",
  3304 => x"808082e3",
  3305 => x"2d848080",
  3306 => x"80932d84",
  3307 => x"8080ecc0",
  3308 => x"51848080",
  3309 => x"82e32d80",
  3310 => x"557483ff",
  3311 => x"e0800c02",
  3312 => x"80c0050d",
  3313 => x"04000000",
  3314 => x"00ffffff",
  3315 => x"ff00ffff",
  3316 => x"ffff00ff",
  3317 => x"ffffff00",
  3318 => x"08200800",
  3319 => x"434d4438",
  3320 => x"5f342072",
  3321 => x"6573706f",
  3322 => x"6e73653a",
  3323 => x"2025640a",
  3324 => x"00000000",
  3325 => x"53444843",
  3326 => x"20496e69",
  3327 => x"7469616c",
  3328 => x"697a6174",
  3329 => x"696f6e20",
  3330 => x"6572726f",
  3331 => x"72210a00",
  3332 => x"434d4435",
  3333 => x"38202564",
  3334 => x"0a202000",
  3335 => x"52656164",
  3336 => x"20636f6d",
  3337 => x"6d616e64",
  3338 => x"20666169",
  3339 => x"6c656420",
  3340 => x"61742025",
  3341 => x"64202825",
  3342 => x"64290a00",
  3343 => x"4641545f",
  3344 => x"46533a20",
  3345 => x"4572726f",
  3346 => x"7220636f",
  3347 => x"756c6420",
  3348 => x"6e6f7420",
  3349 => x"6c6f6164",
  3350 => x"20464154",
  3351 => x"20646574",
  3352 => x"61696c73",
  3353 => x"20282564",
  3354 => x"29210d0a",
  3355 => x"00000000",
  3356 => x"2573203c",
  3357 => x"4449523e",
  3358 => x"0d0a0000",
  3359 => x"2573205b",
  3360 => x"25642062",
  3361 => x"79746573",
  3362 => x"5d0d0a00",
  3363 => x"46415420",
  3364 => x"64657461",
  3365 => x"696c733a",
  3366 => x"0d0a0000",
  3367 => x"46415433",
  3368 => x"32000000",
  3369 => x"46415431",
  3370 => x"36000000",
  3371 => x"20547970",
  3372 => x"65203d25",
  3373 => x"73000000",
  3374 => x"20526f6f",
  3375 => x"74204469",
  3376 => x"72204669",
  3377 => x"72737420",
  3378 => x"436c7573",
  3379 => x"74657220",
  3380 => x"3d202578",
  3381 => x"0d0a0000",
  3382 => x"20464154",
  3383 => x"20426567",
  3384 => x"696e204c",
  3385 => x"4241203d",
  3386 => x"20307825",
  3387 => x"780d0a00",
  3388 => x"20436c75",
  3389 => x"73746572",
  3390 => x"20426567",
  3391 => x"696e204c",
  3392 => x"4241203d",
  3393 => x"20307825",
  3394 => x"780d0a00",
  3395 => x"20536563",
  3396 => x"746f7273",
  3397 => x"20506572",
  3398 => x"20436c75",
  3399 => x"73746572",
  3400 => x"203d2025",
  3401 => x"640d0a00",
  3402 => x"4750494f",
  3403 => x"3020426f",
  3404 => x"6f74206f",
  3405 => x"7074696f",
  3406 => x"6e733a0a",
  3407 => x"00000000",
  3408 => x"30203a20",
  3409 => x"426f6f74",
  3410 => x"2066726f",
  3411 => x"6d205344",
  3412 => x"20636172",
  3413 => x"640a0000",
  3414 => x"31203a20",
  3415 => x"426f6f74",
  3416 => x"2066726f",
  3417 => x"6d204a54",
  3418 => x"41470a00",
  3419 => x"426f6f74",
  3420 => x"696e6720",
  3421 => x"66726f6d",
  3422 => x"20534420",
  3423 => x"63617264",
  3424 => x"0a000000",
  3425 => x"4552524f",
  3426 => x"523a204d",
  3427 => x"65646961",
  3428 => x"20617474",
  3429 => x"61636820",
  3430 => x"6661696c",
  3431 => x"65640a00",
  3432 => x"0a202564",
  3433 => x"20627974",
  3434 => x"65732072",
  3435 => x"6561640a",
  3436 => x"00000000",
  3437 => x"4c697374",
  3438 => x"696e6720",
  3439 => x"64697265",
  3440 => x"63746f72",
  3441 => x"6965732e",
  3442 => x"2e2e0a0a",
  3443 => x"00000000",
  3444 => x"2f000000",
  3445 => x"0a415050",
  3446 => x"2046494c",
  3447 => x"45203e3e",
  3448 => x"20000000",
  3449 => x"72620000",
  3450 => x"0a455252",
  3451 => x"4f523a20",
  3452 => x"52656164",
  3453 => x"2066696c",
  3454 => x"65206661",
  3455 => x"696c6564",
  3456 => x"0a000000",
  3457 => x"426f6f74",
  3458 => x"696e6720",
  3459 => x"66726f6d",
  3460 => x"204a5441",
  3461 => x"472c2077",
  3462 => x"61697469",
  3463 => x"6e672066",
  3464 => x"6f722075",
  3465 => x"706c6f61",
  3466 => x"6465720a",
  3467 => x"00000000",
  3468 => x"454e4400",
  3469 => x"0a0a456e",
  3470 => x"642e2e2e",
  3471 => x"200a0000",
  3472 => x"73687574",
  3473 => x"646f776e",
  3474 => x"2e0a0000",
others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;

		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end rtl;

